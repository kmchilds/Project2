//////////////////////////////////////////////////////////
//														//
//			Written By: Kevin Childs					//
//			Class:		ELEN 249						//
//			Professor:	K. Gunnam & T. Ogunfunmi		//
//			Quarter:	Winter 2016						//
//			Module:		Cosine Generator					//
//			Notes:		Takes in a number between 0 and 1 and gives a cos equiv	//
//														//
//////////////////////////////////////////////////////////


module getCosine2(clk,u1,g0,g1);
input [16:0] u1;
input clk;
output reg [16:0] g0;
output reg [16:0] g1;
wire [16:0] x_g_a;
assign x_g_a = u1[13:0];

wire x_sign, y_sign;
assign x_sign = u1[15];
assign y_sign = u1[14];


reg [16:0] cosLookup[16383:0];


always @(posedge clk)
begin
cosLookup[0] <= 1;
cosLookup[1] <= 0.999999995;
cosLookup[2] <= 0.999999982;
cosLookup[3] <= 0.999999959;
cosLookup[4] <= 0.999999926;
cosLookup[5] <= 0.999999885;
cosLookup[6] <= 0.999999835;
cosLookup[7] <= 0.999999775;
cosLookup[8] <= 0.999999706;
cosLookup[9] <= 0.999999628;
cosLookup[10] <= 0.99999954;
cosLookup[11] <= 0.999999444;
cosLookup[12] <= 0.999999338;
cosLookup[13] <= 0.999999223;
cosLookup[14] <= 0.999999099;
cosLookup[15] <= 0.999998966;
cosLookup[16] <= 0.999998823;
cosLookup[17] <= 0.999998672;
cosLookup[18] <= 0.999998511;
cosLookup[19] <= 0.999998341;
cosLookup[20] <= 0.999998161;
cosLookup[21] <= 0.999997973;
cosLookup[22] <= 0.999997775;
cosLookup[23] <= 0.999997568;
cosLookup[24] <= 0.999997352;
cosLookup[25] <= 0.999997127;
cosLookup[26] <= 0.999996893;
cosLookup[27] <= 0.999996649;
cosLookup[28] <= 0.999996396;
cosLookup[29] <= 0.999996134;
cosLookup[30] <= 0.999995863;
cosLookup[31] <= 0.999995583;
cosLookup[32] <= 0.999995293;
cosLookup[33] <= 0.999994994;
cosLookup[34] <= 0.999994687;
cosLookup[35] <= 0.999994369;
cosLookup[36] <= 0.999994043;
cosLookup[37] <= 0.999993707;
cosLookup[38] <= 0.999993363;
cosLookup[39] <= 0.999993009;
cosLookup[40] <= 0.999992646;
cosLookup[41] <= 0.999992273;
cosLookup[42] <= 0.999991892;
cosLookup[43] <= 0.999991501;
cosLookup[44] <= 0.999991101;
cosLookup[45] <= 0.999990692;
cosLookup[46] <= 0.999990274;
cosLookup[47] <= 0.999989846;
cosLookup[48] <= 0.99998941;
cosLookup[49] <= 0.999988964;
cosLookup[50] <= 0.999988509;
cosLookup[51] <= 0.999988045;
cosLookup[52] <= 0.999987571;
cosLookup[53] <= 0.999987089;
cosLookup[54] <= 0.999986597;
cosLookup[55] <= 0.999986096;
cosLookup[56] <= 0.999985586;
cosLookup[57] <= 0.999985066;
cosLookup[58] <= 0.999984538;
cosLookup[59] <= 0.999984;
cosLookup[60] <= 0.999983453;
cosLookup[61] <= 0.999982897;
cosLookup[62] <= 0.999982331;
cosLookup[63] <= 0.999981757;
cosLookup[64] <= 0.999981173;
cosLookup[65] <= 0.99998058;
cosLookup[66] <= 0.999979978;
cosLookup[67] <= 0.999979367;
cosLookup[68] <= 0.999978746;
cosLookup[69] <= 0.999978116;
cosLookup[70] <= 0.999977477;
cosLookup[71] <= 0.999976829;
cosLookup[72] <= 0.999976172;
cosLookup[73] <= 0.999975506;
cosLookup[74] <= 0.99997483;
cosLookup[75] <= 0.999974145;
cosLookup[76] <= 0.999973451;
cosLookup[77] <= 0.999972748;
cosLookup[78] <= 0.999972035;
cosLookup[79] <= 0.999971314;
cosLookup[80] <= 0.999970583;
cosLookup[81] <= 0.999969843;
cosLookup[82] <= 0.999969094;
cosLookup[83] <= 0.999968335;
cosLookup[84] <= 0.999967568;
cosLookup[85] <= 0.999966791;
cosLookup[86] <= 0.999966005;
cosLookup[87] <= 0.99996521;
cosLookup[88] <= 0.999964405;
cosLookup[89] <= 0.999963592;
cosLookup[90] <= 0.999962769;
cosLookup[91] <= 0.999961937;
cosLookup[92] <= 0.999961096;
cosLookup[93] <= 0.999960246;
cosLookup[94] <= 0.999959386;
cosLookup[95] <= 0.999958517;
cosLookup[96] <= 0.999957639;
cosLookup[97] <= 0.999956752;
cosLookup[98] <= 0.999955856;
cosLookup[99] <= 0.99995495;
cosLookup[100] <= 0.999954036;
cosLookup[101] <= 0.999953112;
cosLookup[102] <= 0.999952179;
cosLookup[103] <= 0.999951237;
cosLookup[104] <= 0.999950285;
cosLookup[105] <= 0.999949325;
cosLookup[106] <= 0.999948355;
cosLookup[107] <= 0.999947376;
cosLookup[108] <= 0.999946387;
cosLookup[109] <= 0.99994539;
cosLookup[110] <= 0.999944383;
cosLookup[111] <= 0.999943368;
cosLookup[112] <= 0.999942343;
cosLookup[113] <= 0.999941308;
cosLookup[114] <= 0.999940265;
cosLookup[115] <= 0.999939213;
cosLookup[116] <= 0.999938151;
cosLookup[117] <= 0.99993708;
cosLookup[118] <= 0.999936;
cosLookup[119] <= 0.99993491;
cosLookup[120] <= 0.999933812;
cosLookup[121] <= 0.999932704;
cosLookup[122] <= 0.999931587;
cosLookup[123] <= 0.999930461;
cosLookup[124] <= 0.999929326;
cosLookup[125] <= 0.999928181;
cosLookup[126] <= 0.999927028;
cosLookup[127] <= 0.999925865;
cosLookup[128] <= 0.999924693;
cosLookup[129] <= 0.999923511;
cosLookup[130] <= 0.999922321;
cosLookup[131] <= 0.999921121;
cosLookup[132] <= 0.999919912;
cosLookup[133] <= 0.999918694;
cosLookup[134] <= 0.999917467;
cosLookup[135] <= 0.999916231;
cosLookup[136] <= 0.999914985;
cosLookup[137] <= 0.99991373;
cosLookup[138] <= 0.999912466;
cosLookup[139] <= 0.999911193;
cosLookup[140] <= 0.999909911;
cosLookup[141] <= 0.999908619;
cosLookup[142] <= 0.999907319;
cosLookup[143] <= 0.999906009;
cosLookup[144] <= 0.999904689;
cosLookup[145] <= 0.999903361;
cosLookup[146] <= 0.999902024;
cosLookup[147] <= 0.999900677;
cosLookup[148] <= 0.999899321;
cosLookup[149] <= 0.999897956;
cosLookup[150] <= 0.999896582;
cosLookup[151] <= 0.999895198;
cosLookup[152] <= 0.999893805;
cosLookup[153] <= 0.999892404;
cosLookup[154] <= 0.999890992;
cosLookup[155] <= 0.999889572;
cosLookup[156] <= 0.999888143;
cosLookup[157] <= 0.999886704;
cosLookup[158] <= 0.999885256;
cosLookup[159] <= 0.999883799;
cosLookup[160] <= 0.999882333;
cosLookup[161] <= 0.999880858;
cosLookup[162] <= 0.999879373;
cosLookup[163] <= 0.999877879;
cosLookup[164] <= 0.999876376;
cosLookup[165] <= 0.999874864;
cosLookup[166] <= 0.999873343;
cosLookup[167] <= 0.999871812;
cosLookup[168] <= 0.999870272;
cosLookup[169] <= 0.999868724;
cosLookup[170] <= 0.999867165;
cosLookup[171] <= 0.999865598;
cosLookup[172] <= 0.999864022;
cosLookup[173] <= 0.999862436;
cosLookup[174] <= 0.999860841;
cosLookup[175] <= 0.999859237;
cosLookup[176] <= 0.999857624;
cosLookup[177] <= 0.999856001;
cosLookup[178] <= 0.999854369;
cosLookup[179] <= 0.999852729;
cosLookup[180] <= 0.999851079;
cosLookup[181] <= 0.999849419;
cosLookup[182] <= 0.999847751;
cosLookup[183] <= 0.999846073;
cosLookup[184] <= 0.999844386;
cosLookup[185] <= 0.99984269;
cosLookup[186] <= 0.999840985;
cosLookup[187] <= 0.999839271;
cosLookup[188] <= 0.999837547;
cosLookup[189] <= 0.999835815;
cosLookup[190] <= 0.999834073;
cosLookup[191] <= 0.999832321;
cosLookup[192] <= 0.999830561;
cosLookup[193] <= 0.999828792;
cosLookup[194] <= 0.999827013;
cosLookup[195] <= 0.999825225;
cosLookup[196] <= 0.999823428;
cosLookup[197] <= 0.999821622;
cosLookup[198] <= 0.999819806;
cosLookup[199] <= 0.999817981;
cosLookup[200] <= 0.999816147;
cosLookup[201] <= 0.999814304;
cosLookup[202] <= 0.999812452;
cosLookup[203] <= 0.999810591;
cosLookup[204] <= 0.99980872;
cosLookup[205] <= 0.99980684;
cosLookup[206] <= 0.999804951;
cosLookup[207] <= 0.999803053;
cosLookup[208] <= 0.999801146;
cosLookup[209] <= 0.999799229;
cosLookup[210] <= 0.999797303;
cosLookup[211] <= 0.999795368;
cosLookup[212] <= 0.999793424;
cosLookup[213] <= 0.999791471;
cosLookup[214] <= 0.999789508;
cosLookup[215] <= 0.999787536;
cosLookup[216] <= 0.999785556;
cosLookup[217] <= 0.999783565;
cosLookup[218] <= 0.999781566;
cosLookup[219] <= 0.999779558;
cosLookup[220] <= 0.99977754;
cosLookup[221] <= 0.999775513;
cosLookup[222] <= 0.999773477;
cosLookup[223] <= 0.999771432;
cosLookup[224] <= 0.999769377;
cosLookup[225] <= 0.999767314;
cosLookup[226] <= 0.999765241;
cosLookup[227] <= 0.999763159;
cosLookup[228] <= 0.999761067;
cosLookup[229] <= 0.999758967;
cosLookup[230] <= 0.999756857;
cosLookup[231] <= 0.999754739;
cosLookup[232] <= 0.999752611;
cosLookup[233] <= 0.999750473;
cosLookup[234] <= 0.999748327;
cosLookup[235] <= 0.999746172;
cosLookup[236] <= 0.999744007;
cosLookup[237] <= 0.999741833;
cosLookup[238] <= 0.99973965;
cosLookup[239] <= 0.999737457;
cosLookup[240] <= 0.999735256;
cosLookup[241] <= 0.999733045;
cosLookup[242] <= 0.999730825;
cosLookup[243] <= 0.999728596;
cosLookup[244] <= 0.999726358;
cosLookup[245] <= 0.999724111;
cosLookup[246] <= 0.999721854;
cosLookup[247] <= 0.999719588;
cosLookup[248] <= 0.999717313;
cosLookup[249] <= 0.999715029;
cosLookup[250] <= 0.999712735;
cosLookup[251] <= 0.999710433;
cosLookup[252] <= 0.999708121;
cosLookup[253] <= 0.9997058;
cosLookup[254] <= 0.99970347;
cosLookup[255] <= 0.99970113;
cosLookup[256] <= 0.999698782;
cosLookup[257] <= 0.999696424;
cosLookup[258] <= 0.999694057;
cosLookup[259] <= 0.999691681;
cosLookup[260] <= 0.999689296;
cosLookup[261] <= 0.999686901;
cosLookup[262] <= 0.999684498;
cosLookup[263] <= 0.999682085;
cosLookup[264] <= 0.999679663;
cosLookup[265] <= 0.999677231;
cosLookup[266] <= 0.999674791;
cosLookup[267] <= 0.999672341;
cosLookup[268] <= 0.999669882;
cosLookup[269] <= 0.999667414;
cosLookup[270] <= 0.999664937;
cosLookup[271] <= 0.999662451;
cosLookup[272] <= 0.999659955;
cosLookup[273] <= 0.99965745;
cosLookup[274] <= 0.999654936;
cosLookup[275] <= 0.999652413;
cosLookup[276] <= 0.999649881;
cosLookup[277] <= 0.999647339;
cosLookup[278] <= 0.999644789;
cosLookup[279] <= 0.999642229;
cosLookup[280] <= 0.99963966;
cosLookup[281] <= 0.999637081;
cosLookup[282] <= 0.999634494;
cosLookup[283] <= 0.999631897;
cosLookup[284] <= 0.999629291;
cosLookup[285] <= 0.999626676;
cosLookup[286] <= 0.999624052;
cosLookup[287] <= 0.999621419;
cosLookup[288] <= 0.999618776;
cosLookup[289] <= 0.999616124;
cosLookup[290] <= 0.999613463;
cosLookup[291] <= 0.999610793;
cosLookup[292] <= 0.999608114;
cosLookup[293] <= 0.999605425;
cosLookup[294] <= 0.999602727;
cosLookup[295] <= 0.99960002;
cosLookup[296] <= 0.999597304;
cosLookup[297] <= 0.999594579;
cosLookup[298] <= 0.999591844;
cosLookup[299] <= 0.999589101;
cosLookup[300] <= 0.999586348;
cosLookup[301] <= 0.999583586;
cosLookup[302] <= 0.999580814;
cosLookup[303] <= 0.999578034;
cosLookup[304] <= 0.999575244;
cosLookup[305] <= 0.999572445;
cosLookup[306] <= 0.999569637;
cosLookup[307] <= 0.99956682;
cosLookup[308] <= 0.999563994;
cosLookup[309] <= 0.999561158;
cosLookup[310] <= 0.999558313;
cosLookup[311] <= 0.999555459;
cosLookup[312] <= 0.999552596;
cosLookup[313] <= 0.999549724;
cosLookup[314] <= 0.999546842;
cosLookup[315] <= 0.999543952;
cosLookup[316] <= 0.999541052;
cosLookup[317] <= 0.999538143;
cosLookup[318] <= 0.999535224;
cosLookup[319] <= 0.999532297;
cosLookup[320] <= 0.99952936;
cosLookup[321] <= 0.999526414;
cosLookup[322] <= 0.999523459;
cosLookup[323] <= 0.999520495;
cosLookup[324] <= 0.999517521;
cosLookup[325] <= 0.999514539;
cosLookup[326] <= 0.999511547;
cosLookup[327] <= 0.999508546;
cosLookup[328] <= 0.999505536;
cosLookup[329] <= 0.999502517;
cosLookup[330] <= 0.999499488;
cosLookup[331] <= 0.99949645;
cosLookup[332] <= 0.999493403;
cosLookup[333] <= 0.999490347;
cosLookup[334] <= 0.999487282;
cosLookup[335] <= 0.999484207;
cosLookup[336] <= 0.999481124;
cosLookup[337] <= 0.999478031;
cosLookup[338] <= 0.999474929;
cosLookup[339] <= 0.999471817;
cosLookup[340] <= 0.999468697;
cosLookup[341] <= 0.999465567;
cosLookup[342] <= 0.999462429;
cosLookup[343] <= 0.999459281;
cosLookup[344] <= 0.999456123;
cosLookup[345] <= 0.999452957;
cosLookup[346] <= 0.999449781;
cosLookup[347] <= 0.999446597;
cosLookup[348] <= 0.999443403;
cosLookup[349] <= 0.9994402;
cosLookup[350] <= 0.999436987;
cosLookup[351] <= 0.999433766;
cosLookup[352] <= 0.999430535;
cosLookup[353] <= 0.999427295;
cosLookup[354] <= 0.999424046;
cosLookup[355] <= 0.999420788;
cosLookup[356] <= 0.99941752;
cosLookup[357] <= 0.999414244;
cosLookup[358] <= 0.999410958;
cosLookup[359] <= 0.999407663;
cosLookup[360] <= 0.999404359;
cosLookup[361] <= 0.999401045;
cosLookup[362] <= 0.999397723;
cosLookup[363] <= 0.999394391;
cosLookup[364] <= 0.99939105;
cosLookup[365] <= 0.9993877;
cosLookup[366] <= 0.999384341;
cosLookup[367] <= 0.999380972;
cosLookup[368] <= 0.999377594;
cosLookup[369] <= 0.999374208;
cosLookup[370] <= 0.999370811;
cosLookup[371] <= 0.999367406;
cosLookup[372] <= 0.999363992;
cosLookup[373] <= 0.999360568;
cosLookup[374] <= 0.999357135;
cosLookup[375] <= 0.999353693;
cosLookup[376] <= 0.999350242;
cosLookup[377] <= 0.999346782;
cosLookup[378] <= 0.999343312;
cosLookup[379] <= 0.999339833;
cosLookup[380] <= 0.999336345;
cosLookup[381] <= 0.999332848;
cosLookup[382] <= 0.999329342;
cosLookup[383] <= 0.999325827;
cosLookup[384] <= 0.999322302;
cosLookup[385] <= 0.999318768;
cosLookup[386] <= 0.999315225;
cosLookup[387] <= 0.999311673;
cosLookup[388] <= 0.999308111;
cosLookup[389] <= 0.999304541;
cosLookup[390] <= 0.999300961;
cosLookup[391] <= 0.999297372;
cosLookup[392] <= 0.999293774;
cosLookup[393] <= 0.999290166;
cosLookup[394] <= 0.99928655;
cosLookup[395] <= 0.999282924;
cosLookup[396] <= 0.999279289;
cosLookup[397] <= 0.999275645;
cosLookup[398] <= 0.999271992;
cosLookup[399] <= 0.999268329;
cosLookup[400] <= 0.999264658;
cosLookup[401] <= 0.999260977;
cosLookup[402] <= 0.999257287;
cosLookup[403] <= 0.999253587;
cosLookup[404] <= 0.999249879;
cosLookup[405] <= 0.999246161;
cosLookup[406] <= 0.999242435;
cosLookup[407] <= 0.999238699;
cosLookup[408] <= 0.999234953;
cosLookup[409] <= 0.999231199;
cosLookup[410] <= 0.999227436;
cosLookup[411] <= 0.999223663;
cosLookup[412] <= 0.999219881;
cosLookup[413] <= 0.99921609;
cosLookup[414] <= 0.99921229;
cosLookup[415] <= 0.99920848;
cosLookup[416] <= 0.999204662;
cosLookup[417] <= 0.999200834;
cosLookup[418] <= 0.999196997;
cosLookup[419] <= 0.999193151;
cosLookup[420] <= 0.999189295;
cosLookup[421] <= 0.999185431;
cosLookup[422] <= 0.999181557;
cosLookup[423] <= 0.999177674;
cosLookup[424] <= 0.999173782;
cosLookup[425] <= 0.99916988;
cosLookup[426] <= 0.99916597;
cosLookup[427] <= 0.99916205;
cosLookup[428] <= 0.999158121;
cosLookup[429] <= 0.999154183;
cosLookup[430] <= 0.999150236;
cosLookup[431] <= 0.99914628;
cosLookup[432] <= 0.999142314;
cosLookup[433] <= 0.999138339;
cosLookup[434] <= 0.999134355;
cosLookup[435] <= 0.999130362;
cosLookup[436] <= 0.99912636;
cosLookup[437] <= 0.999122348;
cosLookup[438] <= 0.999118328;
cosLookup[439] <= 0.999114298;
cosLookup[440] <= 0.999110259;
cosLookup[441] <= 0.99910621;
cosLookup[442] <= 0.999102153;
cosLookup[443] <= 0.999098086;
cosLookup[444] <= 0.99909401;
cosLookup[445] <= 0.999089925;
cosLookup[446] <= 0.999085831;
cosLookup[447] <= 0.999081728;
cosLookup[448] <= 0.999077615;
cosLookup[449] <= 0.999073493;
cosLookup[450] <= 0.999069362;
cosLookup[451] <= 0.999065222;
cosLookup[452] <= 0.999061073;
cosLookup[453] <= 0.999056915;
cosLookup[454] <= 0.999052747;
cosLookup[455] <= 0.99904857;
cosLookup[456] <= 0.999044384;
cosLookup[457] <= 0.999040189;
cosLookup[458] <= 0.999035984;
cosLookup[459] <= 0.999031771;
cosLookup[460] <= 0.999027548;
cosLookup[461] <= 0.999023316;
cosLookup[462] <= 0.999019075;
cosLookup[463] <= 0.999014825;
cosLookup[464] <= 0.999010565;
cosLookup[465] <= 0.999006296;
cosLookup[466] <= 0.999002019;
cosLookup[467] <= 0.998997731;
cosLookup[468] <= 0.998993435;
cosLookup[469] <= 0.99898913;
cosLookup[470] <= 0.998984815;
cosLookup[471] <= 0.998980491;
cosLookup[472] <= 0.998976158;
cosLookup[473] <= 0.998971816;
cosLookup[474] <= 0.998967465;
cosLookup[475] <= 0.998963104;
cosLookup[476] <= 0.998958735;
cosLookup[477] <= 0.998954356;
cosLookup[478] <= 0.998949968;
cosLookup[479] <= 0.99894557;
cosLookup[480] <= 0.998941164;
cosLookup[481] <= 0.998936748;
cosLookup[482] <= 0.998932324;
cosLookup[483] <= 0.99892789;
cosLookup[484] <= 0.998923446;
cosLookup[485] <= 0.998918994;
cosLookup[486] <= 0.998914532;
cosLookup[487] <= 0.998910062;
cosLookup[488] <= 0.998905582;
cosLookup[489] <= 0.998901093;
cosLookup[490] <= 0.998896594;
cosLookup[491] <= 0.998892087;
cosLookup[492] <= 0.99888757;
cosLookup[493] <= 0.998883045;
cosLookup[494] <= 0.998878509;
cosLookup[495] <= 0.998873965;
cosLookup[496] <= 0.998869412;
cosLookup[497] <= 0.998864849;
cosLookup[498] <= 0.998860278;
cosLookup[499] <= 0.998855697;
cosLookup[500] <= 0.998851107;
cosLookup[501] <= 0.998846507;
cosLookup[502] <= 0.998841899;
cosLookup[503] <= 0.998837281;
cosLookup[504] <= 0.998832654;
cosLookup[505] <= 0.998828018;
cosLookup[506] <= 0.998823373;
cosLookup[507] <= 0.998818719;
cosLookup[508] <= 0.998814055;
cosLookup[509] <= 0.998809382;
cosLookup[510] <= 0.998804701;
cosLookup[511] <= 0.998800009;
cosLookup[512] <= 0.998795309;
cosLookup[513] <= 0.9987906;
cosLookup[514] <= 0.998785881;
cosLookup[515] <= 0.998781153;
cosLookup[516] <= 0.998776416;
cosLookup[517] <= 0.99877167;
cosLookup[518] <= 0.998766915;
cosLookup[519] <= 0.99876215;
cosLookup[520] <= 0.998757376;
cosLookup[521] <= 0.998752593;
cosLookup[522] <= 0.998747801;
cosLookup[523] <= 0.998743;
cosLookup[524] <= 0.99873819;
cosLookup[525] <= 0.99873337;
cosLookup[526] <= 0.998728541;
cosLookup[527] <= 0.998723703;
cosLookup[528] <= 0.998718856;
cosLookup[529] <= 0.998714;
cosLookup[530] <= 0.998709134;
cosLookup[531] <= 0.998704259;
cosLookup[532] <= 0.998699375;
cosLookup[533] <= 0.998694482;
cosLookup[534] <= 0.99868958;
cosLookup[535] <= 0.998684668;
cosLookup[536] <= 0.998679748;
cosLookup[537] <= 0.998674818;
cosLookup[538] <= 0.998669879;
cosLookup[539] <= 0.998664931;
cosLookup[540] <= 0.998659973;
cosLookup[541] <= 0.998655007;
cosLookup[542] <= 0.998650031;
cosLookup[543] <= 0.998645046;
cosLookup[544] <= 0.998640052;
cosLookup[545] <= 0.998635049;
cosLookup[546] <= 0.998630037;
cosLookup[547] <= 0.998625015;
cosLookup[548] <= 0.998619984;
cosLookup[549] <= 0.998614944;
cosLookup[550] <= 0.998609895;
cosLookup[551] <= 0.998604837;
cosLookup[552] <= 0.998599769;
cosLookup[553] <= 0.998594692;
cosLookup[554] <= 0.998589606;
cosLookup[555] <= 0.998584511;
cosLookup[556] <= 0.998579407;
cosLookup[557] <= 0.998574294;
cosLookup[558] <= 0.998569171;
cosLookup[559] <= 0.998564039;
cosLookup[560] <= 0.998558898;
cosLookup[561] <= 0.998553748;
cosLookup[562] <= 0.998548589;
cosLookup[563] <= 0.99854342;
cosLookup[564] <= 0.998538243;
cosLookup[565] <= 0.998533056;
cosLookup[566] <= 0.99852786;
cosLookup[567] <= 0.998522655;
cosLookup[568] <= 0.99851744;
cosLookup[569] <= 0.998512217;
cosLookup[570] <= 0.998506984;
cosLookup[571] <= 0.998501742;
cosLookup[572] <= 0.998496491;
cosLookup[573] <= 0.99849123;
cosLookup[574] <= 0.998485961;
cosLookup[575] <= 0.998480682;
cosLookup[576] <= 0.998475395;
cosLookup[577] <= 0.998470098;
cosLookup[578] <= 0.998464791;
cosLookup[579] <= 0.998459476;
cosLookup[580] <= 0.998454151;
cosLookup[581] <= 0.998448818;
cosLookup[582] <= 0.998443475;
cosLookup[583] <= 0.998438123;
cosLookup[584] <= 0.998432761;
cosLookup[585] <= 0.998427391;
cosLookup[586] <= 0.998422011;
cosLookup[587] <= 0.998416623;
cosLookup[588] <= 0.998411225;
cosLookup[589] <= 0.998405817;
cosLookup[590] <= 0.998400401;
cosLookup[591] <= 0.998394976;
cosLookup[592] <= 0.998389541;
cosLookup[593] <= 0.998384097;
cosLookup[594] <= 0.998378644;
cosLookup[595] <= 0.998373182;
cosLookup[596] <= 0.99836771;
cosLookup[597] <= 0.99836223;
cosLookup[598] <= 0.99835674;
cosLookup[599] <= 0.998351241;
cosLookup[600] <= 0.998345733;
cosLookup[601] <= 0.998340216;
cosLookup[602] <= 0.998334689;
cosLookup[603] <= 0.998329154;
cosLookup[604] <= 0.998323609;
cosLookup[605] <= 0.998318055;
cosLookup[606] <= 0.998312492;
cosLookup[607] <= 0.998306919;
cosLookup[608] <= 0.998301338;
cosLookup[609] <= 0.998295747;
cosLookup[610] <= 0.998290147;
cosLookup[611] <= 0.998284538;
cosLookup[612] <= 0.99827892;
cosLookup[613] <= 0.998273292;
cosLookup[614] <= 0.998267656;
cosLookup[615] <= 0.99826201;
cosLookup[616] <= 0.998256355;
cosLookup[617] <= 0.998250691;
cosLookup[618] <= 0.998245018;
cosLookup[619] <= 0.998239335;
cosLookup[620] <= 0.998233643;
cosLookup[621] <= 0.998227943;
cosLookup[622] <= 0.998222233;
cosLookup[623] <= 0.998216513;
cosLookup[624] <= 0.998210785;
cosLookup[625] <= 0.998205047;
cosLookup[626] <= 0.998199301;
cosLookup[627] <= 0.998193545;
cosLookup[628] <= 0.99818778;
cosLookup[629] <= 0.998182006;
cosLookup[630] <= 0.998176222;
cosLookup[631] <= 0.99817043;
cosLookup[632] <= 0.998164628;
cosLookup[633] <= 0.998158817;
cosLookup[634] <= 0.998152997;
cosLookup[635] <= 0.998147167;
cosLookup[636] <= 0.998141329;
cosLookup[637] <= 0.998135481;
cosLookup[638] <= 0.998129624;
cosLookup[639] <= 0.998123758;
cosLookup[640] <= 0.998117883;
cosLookup[641] <= 0.998111999;
cosLookup[642] <= 0.998106105;
cosLookup[643] <= 0.998100203;
cosLookup[644] <= 0.998094291;
cosLookup[645] <= 0.99808837;
cosLookup[646] <= 0.998082439;
cosLookup[647] <= 0.9980765;
cosLookup[648] <= 0.998070551;
cosLookup[649] <= 0.998064594;
cosLookup[650] <= 0.998058627;
cosLookup[651] <= 0.998052651;
cosLookup[652] <= 0.998046665;
cosLookup[653] <= 0.998040671;
cosLookup[654] <= 0.998034667;
cosLookup[655] <= 0.998028654;
cosLookup[656] <= 0.998022632;
cosLookup[657] <= 0.998016601;
cosLookup[658] <= 0.998010561;
cosLookup[659] <= 0.998004511;
cosLookup[660] <= 0.997998453;
cosLookup[661] <= 0.997992385;
cosLookup[662] <= 0.997986308;
cosLookup[663] <= 0.997980222;
cosLookup[664] <= 0.997974126;
cosLookup[665] <= 0.997968022;
cosLookup[666] <= 0.997961908;
cosLookup[667] <= 0.997955785;
cosLookup[668] <= 0.997949653;
cosLookup[669] <= 0.997943512;
cosLookup[670] <= 0.997937361;
cosLookup[671] <= 0.997931202;
cosLookup[672] <= 0.997925033;
cosLookup[673] <= 0.997918855;
cosLookup[674] <= 0.997912668;
cosLookup[675] <= 0.997906472;
cosLookup[676] <= 0.997900266;
cosLookup[677] <= 0.997894052;
cosLookup[678] <= 0.997887828;
cosLookup[679] <= 0.997881595;
cosLookup[680] <= 0.997875353;
cosLookup[681] <= 0.997869101;
cosLookup[682] <= 0.997862841;
cosLookup[683] <= 0.997856571;
cosLookup[684] <= 0.997850292;
cosLookup[685] <= 0.997844004;
cosLookup[686] <= 0.997837707;
cosLookup[687] <= 0.997831401;
cosLookup[688] <= 0.997825085;
cosLookup[689] <= 0.99781876;
cosLookup[690] <= 0.997812426;
cosLookup[691] <= 0.997806083;
cosLookup[692] <= 0.997799731;
cosLookup[693] <= 0.99779337;
cosLookup[694] <= 0.997786999;
cosLookup[695] <= 0.997780619;
cosLookup[696] <= 0.99777423;
cosLookup[697] <= 0.997767832;
cosLookup[698] <= 0.997761425;
cosLookup[699] <= 0.997755009;
cosLookup[700] <= 0.997748583;
cosLookup[701] <= 0.997742148;
cosLookup[702] <= 0.997735704;
cosLookup[703] <= 0.997729251;
cosLookup[704] <= 0.997722789;
cosLookup[705] <= 0.997716317;
cosLookup[706] <= 0.997709837;
cosLookup[707] <= 0.997703347;
cosLookup[708] <= 0.997696848;
cosLookup[709] <= 0.99769034;
cosLookup[710] <= 0.997683822;
cosLookup[711] <= 0.997677296;
cosLookup[712] <= 0.99767076;
cosLookup[713] <= 0.997664215;
cosLookup[714] <= 0.997657661;
cosLookup[715] <= 0.997651098;
cosLookup[716] <= 0.997644526;
cosLookup[717] <= 0.997637944;
cosLookup[718] <= 0.997631353;
cosLookup[719] <= 0.997624754;
cosLookup[720] <= 0.997618145;
cosLookup[721] <= 0.997611526;
cosLookup[722] <= 0.997604899;
cosLookup[723] <= 0.997598262;
cosLookup[724] <= 0.997591617;
cosLookup[725] <= 0.997584962;
cosLookup[726] <= 0.997578298;
cosLookup[727] <= 0.997571624;
cosLookup[728] <= 0.997564942;
cosLookup[729] <= 0.99755825;
cosLookup[730] <= 0.99755155;
cosLookup[731] <= 0.99754484;
cosLookup[732] <= 0.997538121;
cosLookup[733] <= 0.997531392;
cosLookup[734] <= 0.997524655;
cosLookup[735] <= 0.997517908;
cosLookup[736] <= 0.997511152;
cosLookup[737] <= 0.997504388;
cosLookup[738] <= 0.997497613;
cosLookup[739] <= 0.99749083;
cosLookup[740] <= 0.997484038;
cosLookup[741] <= 0.997477236;
cosLookup[742] <= 0.997470425;
cosLookup[743] <= 0.997463605;
cosLookup[744] <= 0.997456776;
cosLookup[745] <= 0.997449938;
cosLookup[746] <= 0.99744309;
cosLookup[747] <= 0.997436234;
cosLookup[748] <= 0.997429368;
cosLookup[749] <= 0.997422493;
cosLookup[750] <= 0.997415609;
cosLookup[751] <= 0.997408715;
cosLookup[752] <= 0.997401813;
cosLookup[753] <= 0.997394901;
cosLookup[754] <= 0.99738798;
cosLookup[755] <= 0.99738105;
cosLookup[756] <= 0.997374111;
cosLookup[757] <= 0.997367163;
cosLookup[758] <= 0.997360205;
cosLookup[759] <= 0.997353239;
cosLookup[760] <= 0.997346263;
cosLookup[761] <= 0.997339278;
cosLookup[762] <= 0.997332284;
cosLookup[763] <= 0.99732528;
cosLookup[764] <= 0.997318268;
cosLookup[765] <= 0.997311246;
cosLookup[766] <= 0.997304215;
cosLookup[767] <= 0.997297175;
cosLookup[768] <= 0.997290126;
cosLookup[769] <= 0.997283068;
cosLookup[770] <= 0.997276;
cosLookup[771] <= 0.997268923;
cosLookup[772] <= 0.997261838;
cosLookup[773] <= 0.997254743;
cosLookup[774] <= 0.997247638;
cosLookup[775] <= 0.997240525;
cosLookup[776] <= 0.997233402;
cosLookup[777] <= 0.997226271;
cosLookup[778] <= 0.99721913;
cosLookup[779] <= 0.99721198;
cosLookup[780] <= 0.997204821;
cosLookup[781] <= 0.997197652;
cosLookup[782] <= 0.997190475;
cosLookup[783] <= 0.997183288;
cosLookup[784] <= 0.997176092;
cosLookup[785] <= 0.997168887;
cosLookup[786] <= 0.997161673;
cosLookup[787] <= 0.99715445;
cosLookup[788] <= 0.997147217;
cosLookup[789] <= 0.997139975;
cosLookup[790] <= 0.997132724;
cosLookup[791] <= 0.997125464;
cosLookup[792] <= 0.997118195;
cosLookup[793] <= 0.997110917;
cosLookup[794] <= 0.997103629;
cosLookup[795] <= 0.997096333;
cosLookup[796] <= 0.997089027;
cosLookup[797] <= 0.997081712;
cosLookup[798] <= 0.997074388;
cosLookup[799] <= 0.997067054;
cosLookup[800] <= 0.997059712;
cosLookup[801] <= 0.99705236;
cosLookup[802] <= 0.997044999;
cosLookup[803] <= 0.997037629;
cosLookup[804] <= 0.99703025;
cosLookup[805] <= 0.997022861;
cosLookup[806] <= 0.997015464;
cosLookup[807] <= 0.997008057;
cosLookup[808] <= 0.997000641;
cosLookup[809] <= 0.996993216;
cosLookup[810] <= 0.996985782;
cosLookup[811] <= 0.996978339;
cosLookup[812] <= 0.996970886;
cosLookup[813] <= 0.996963425;
cosLookup[814] <= 0.996955954;
cosLookup[815] <= 0.996948474;
cosLookup[816] <= 0.996940985;
cosLookup[817] <= 0.996933486;
cosLookup[818] <= 0.996925979;
cosLookup[819] <= 0.996918462;
cosLookup[820] <= 0.996910936;
cosLookup[821] <= 0.996903401;
cosLookup[822] <= 0.996895857;
cosLookup[823] <= 0.996888304;
cosLookup[824] <= 0.996880741;
cosLookup[825] <= 0.99687317;
cosLookup[826] <= 0.996865589;
cosLookup[827] <= 0.996857999;
cosLookup[828] <= 0.9968504;
cosLookup[829] <= 0.996842791;
cosLookup[830] <= 0.996835174;
cosLookup[831] <= 0.996827547;
cosLookup[832] <= 0.996819911;
cosLookup[833] <= 0.996812266;
cosLookup[834] <= 0.996804612;
cosLookup[835] <= 0.996796949;
cosLookup[836] <= 0.996789276;
cosLookup[837] <= 0.996781595;
cosLookup[838] <= 0.996773904;
cosLookup[839] <= 0.996766204;
cosLookup[840] <= 0.996758495;
cosLookup[841] <= 0.996750777;
cosLookup[842] <= 0.996743049;
cosLookup[843] <= 0.996735313;
cosLookup[844] <= 0.996727567;
cosLookup[845] <= 0.996719812;
cosLookup[846] <= 0.996712048;
cosLookup[847] <= 0.996704275;
cosLookup[848] <= 0.996696492;
cosLookup[849] <= 0.996688701;
cosLookup[850] <= 0.9966809;
cosLookup[851] <= 0.99667309;
cosLookup[852] <= 0.996665271;
cosLookup[853] <= 0.996657443;
cosLookup[854] <= 0.996649605;
cosLookup[855] <= 0.996641759;
cosLookup[856] <= 0.996633903;
cosLookup[857] <= 0.996626038;
cosLookup[858] <= 0.996618164;
cosLookup[859] <= 0.996610281;
cosLookup[860] <= 0.996602389;
cosLookup[861] <= 0.996594487;
cosLookup[862] <= 0.996586576;
cosLookup[863] <= 0.996578656;
cosLookup[864] <= 0.996570727;
cosLookup[865] <= 0.996562789;
cosLookup[866] <= 0.996554842;
cosLookup[867] <= 0.996546885;
cosLookup[868] <= 0.99653892;
cosLookup[869] <= 0.996530945;
cosLookup[870] <= 0.996522961;
cosLookup[871] <= 0.996514968;
cosLookup[872] <= 0.996506966;
cosLookup[873] <= 0.996498954;
cosLookup[874] <= 0.996490933;
cosLookup[875] <= 0.996482904;
cosLookup[876] <= 0.996474865;
cosLookup[877] <= 0.996466817;
cosLookup[878] <= 0.996458759;
cosLookup[879] <= 0.996450693;
cosLookup[880] <= 0.996442617;
cosLookup[881] <= 0.996434533;
cosLookup[882] <= 0.996426439;
cosLookup[883] <= 0.996418336;
cosLookup[884] <= 0.996410223;
cosLookup[885] <= 0.996402102;
cosLookup[886] <= 0.996393972;
cosLookup[887] <= 0.996385832;
cosLookup[888] <= 0.996377683;
cosLookup[889] <= 0.996369525;
cosLookup[890] <= 0.996361358;
cosLookup[891] <= 0.996353181;
cosLookup[892] <= 0.996344996;
cosLookup[893] <= 0.996336801;
cosLookup[894] <= 0.996328597;
cosLookup[895] <= 0.996320384;
cosLookup[896] <= 0.996312162;
cosLookup[897] <= 0.996303931;
cosLookup[898] <= 0.996295691;
cosLookup[899] <= 0.996287441;
cosLookup[900] <= 0.996279182;
cosLookup[901] <= 0.996270914;
cosLookup[902] <= 0.996262637;
cosLookup[903] <= 0.996254351;
cosLookup[904] <= 0.996246055;
cosLookup[905] <= 0.996237751;
cosLookup[906] <= 0.996229437;
cosLookup[907] <= 0.996221114;
cosLookup[908] <= 0.996212782;
cosLookup[909] <= 0.996204441;
cosLookup[910] <= 0.996196091;
cosLookup[911] <= 0.996187731;
cosLookup[912] <= 0.996179363;
cosLookup[913] <= 0.996170985;
cosLookup[914] <= 0.996162598;
cosLookup[915] <= 0.996154202;
cosLookup[916] <= 0.996145796;
cosLookup[917] <= 0.996137382;
cosLookup[918] <= 0.996128958;
cosLookup[919] <= 0.996120525;
cosLookup[920] <= 0.996112083;
cosLookup[921] <= 0.996103632;
cosLookup[922] <= 0.996095172;
cosLookup[923] <= 0.996086703;
cosLookup[924] <= 0.996078224;
cosLookup[925] <= 0.996069736;
cosLookup[926] <= 0.99606124;
cosLookup[927] <= 0.996052734;
cosLookup[928] <= 0.996044218;
cosLookup[929] <= 0.996035694;
cosLookup[930] <= 0.996027161;
cosLookup[931] <= 0.996018618;
cosLookup[932] <= 0.996010066;
cosLookup[933] <= 0.996001505;
cosLookup[934] <= 0.995992935;
cosLookup[935] <= 0.995984356;
cosLookup[936] <= 0.995975767;
cosLookup[937] <= 0.99596717;
cosLookup[938] <= 0.995958563;
cosLookup[939] <= 0.995949947;
cosLookup[940] <= 0.995941322;
cosLookup[941] <= 0.995932688;
cosLookup[942] <= 0.995924044;
cosLookup[943] <= 0.995915392;
cosLookup[944] <= 0.99590673;
cosLookup[945] <= 0.995898059;
cosLookup[946] <= 0.995889379;
cosLookup[947] <= 0.99588069;
cosLookup[948] <= 0.995871992;
cosLookup[949] <= 0.995863284;
cosLookup[950] <= 0.995854568;
cosLookup[951] <= 0.995845842;
cosLookup[952] <= 0.995837107;
cosLookup[953] <= 0.995828363;
cosLookup[954] <= 0.99581961;
cosLookup[955] <= 0.995810847;
cosLookup[956] <= 0.995802076;
cosLookup[957] <= 0.995793295;
cosLookup[958] <= 0.995784505;
cosLookup[959] <= 0.995775706;
cosLookup[960] <= 0.995766898;
cosLookup[961] <= 0.995758081;
cosLookup[962] <= 0.995749254;
cosLookup[963] <= 0.995740419;
cosLookup[964] <= 0.995731574;
cosLookup[965] <= 0.99572272;
cosLookup[966] <= 0.995713857;
cosLookup[967] <= 0.995704985;
cosLookup[968] <= 0.995696103;
cosLookup[969] <= 0.995687213;
cosLookup[970] <= 0.995678313;
cosLookup[971] <= 0.995669404;
cosLookup[972] <= 0.995660486;
cosLookup[973] <= 0.995651559;
cosLookup[974] <= 0.995642623;
cosLookup[975] <= 0.995633677;
cosLookup[976] <= 0.995624723;
cosLookup[977] <= 0.995615759;
cosLookup[978] <= 0.995606786;
cosLookup[979] <= 0.995597804;
cosLookup[980] <= 0.995588813;
cosLookup[981] <= 0.995579812;
cosLookup[982] <= 0.995570803;
cosLookup[983] <= 0.995561784;
cosLookup[984] <= 0.995552756;
cosLookup[985] <= 0.995543719;
cosLookup[986] <= 0.995534673;
cosLookup[987] <= 0.995525618;
cosLookup[988] <= 0.995516553;
cosLookup[989] <= 0.99550748;
cosLookup[990] <= 0.995498397;
cosLookup[991] <= 0.995489305;
cosLookup[992] <= 0.995480204;
cosLookup[993] <= 0.995471094;
cosLookup[994] <= 0.995461975;
cosLookup[995] <= 0.995452846;
cosLookup[996] <= 0.995443708;
cosLookup[997] <= 0.995434562;
cosLookup[998] <= 0.995425406;
cosLookup[999] <= 0.995416241;
cosLookup[1000] <= 0.995407066;
cosLookup[1001] <= 0.995397883;
cosLookup[1002] <= 0.99538869;
cosLookup[1003] <= 0.995379489;
cosLookup[1004] <= 0.995370278;
cosLookup[1005] <= 0.995361058;
cosLookup[1006] <= 0.995351829;
cosLookup[1007] <= 0.99534259;
cosLookup[1008] <= 0.995333343;
cosLookup[1009] <= 0.995324086;
cosLookup[1010] <= 0.995314821;
cosLookup[1011] <= 0.995305546;
cosLookup[1012] <= 0.995296262;
cosLookup[1013] <= 0.995286968;
cosLookup[1014] <= 0.995277666;
cosLookup[1015] <= 0.995268355;
cosLookup[1016] <= 0.995259034;
cosLookup[1017] <= 0.995249704;
cosLookup[1018] <= 0.995240365;
cosLookup[1019] <= 0.995231017;
cosLookup[1020] <= 0.99522166;
cosLookup[1021] <= 0.995212293;
cosLookup[1022] <= 0.995202918;
cosLookup[1023] <= 0.995193533;
cosLookup[1024] <= 0.995184139;
cosLookup[1025] <= 0.995174736;
cosLookup[1026] <= 0.995165324;
cosLookup[1027] <= 0.995155903;
cosLookup[1028] <= 0.995146472;
cosLookup[1029] <= 0.995137033;
cosLookup[1030] <= 0.995127584;
cosLookup[1031] <= 0.995118126;
cosLookup[1032] <= 0.995108659;
cosLookup[1033] <= 0.995099183;
cosLookup[1034] <= 0.995089698;
cosLookup[1035] <= 0.995080203;
cosLookup[1036] <= 0.9950707;
cosLookup[1037] <= 0.995061187;
cosLookup[1038] <= 0.995051665;
cosLookup[1039] <= 0.995042134;
cosLookup[1040] <= 0.995032594;
cosLookup[1041] <= 0.995023044;
cosLookup[1042] <= 0.995013486;
cosLookup[1043] <= 0.995003918;
cosLookup[1044] <= 0.994994341;
cosLookup[1045] <= 0.994984755;
cosLookup[1046] <= 0.99497516;
cosLookup[1047] <= 0.994965556;
cosLookup[1048] <= 0.994955943;
cosLookup[1049] <= 0.99494632;
cosLookup[1050] <= 0.994936688;
cosLookup[1051] <= 0.994927048;
cosLookup[1052] <= 0.994917398;
cosLookup[1053] <= 0.994907738;
cosLookup[1054] <= 0.99489807;
cosLookup[1055] <= 0.994888393;
cosLookup[1056] <= 0.994878706;
cosLookup[1057] <= 0.99486901;
cosLookup[1058] <= 0.994859306;
cosLookup[1059] <= 0.994849592;
cosLookup[1060] <= 0.994839868;
cosLookup[1061] <= 0.994830136;
cosLookup[1062] <= 0.994820395;
cosLookup[1063] <= 0.994810644;
cosLookup[1064] <= 0.994800884;
cosLookup[1065] <= 0.994791116;
cosLookup[1066] <= 0.994781338;
cosLookup[1067] <= 0.99477155;
cosLookup[1068] <= 0.994761754;
cosLookup[1069] <= 0.994751949;
cosLookup[1070] <= 0.994742134;
cosLookup[1071] <= 0.99473231;
cosLookup[1072] <= 0.994722477;
cosLookup[1073] <= 0.994712635;
cosLookup[1074] <= 0.994702784;
cosLookup[1075] <= 0.994692924;
cosLookup[1076] <= 0.994683054;
cosLookup[1077] <= 0.994673176;
cosLookup[1078] <= 0.994663288;
cosLookup[1079] <= 0.994653391;
cosLookup[1080] <= 0.994643485;
cosLookup[1081] <= 0.99463357;
cosLookup[1082] <= 0.994623646;
cosLookup[1083] <= 0.994613712;
cosLookup[1084] <= 0.99460377;
cosLookup[1085] <= 0.994593818;
cosLookup[1086] <= 0.994583857;
cosLookup[1087] <= 0.994573887;
cosLookup[1088] <= 0.994563908;
cosLookup[1089] <= 0.994553919;
cosLookup[1090] <= 0.994543922;
cosLookup[1091] <= 0.994533915;
cosLookup[1092] <= 0.9945239;
cosLookup[1093] <= 0.994513875;
cosLookup[1094] <= 0.994503841;
cosLookup[1095] <= 0.994493798;
cosLookup[1096] <= 0.994483745;
cosLookup[1097] <= 0.994473684;
cosLookup[1098] <= 0.994463613;
cosLookup[1099] <= 0.994453533;
cosLookup[1100] <= 0.994443444;
cosLookup[1101] <= 0.994433346;
cosLookup[1102] <= 0.994423239;
cosLookup[1103] <= 0.994413123;
cosLookup[1104] <= 0.994402997;
cosLookup[1105] <= 0.994392863;
cosLookup[1106] <= 0.994382719;
cosLookup[1107] <= 0.994372566;
cosLookup[1108] <= 0.994362404;
cosLookup[1109] <= 0.994352233;
cosLookup[1110] <= 0.994342053;
cosLookup[1111] <= 0.994331863;
cosLookup[1112] <= 0.994321665;
cosLookup[1113] <= 0.994311457;
cosLookup[1114] <= 0.99430124;
cosLookup[1115] <= 0.994291014;
cosLookup[1116] <= 0.994280779;
cosLookup[1117] <= 0.994270535;
cosLookup[1118] <= 0.994260281;
cosLookup[1119] <= 0.994250019;
cosLookup[1120] <= 0.994239747;
cosLookup[1121] <= 0.994229466;
cosLookup[1122] <= 0.994219176;
cosLookup[1123] <= 0.994208877;
cosLookup[1124] <= 0.994198569;
cosLookup[1125] <= 0.994188251;
cosLookup[1126] <= 0.994177925;
cosLookup[1127] <= 0.994167589;
cosLookup[1128] <= 0.994157244;
cosLookup[1129] <= 0.99414689;
cosLookup[1130] <= 0.994136527;
cosLookup[1131] <= 0.994126155;
cosLookup[1132] <= 0.994115774;
cosLookup[1133] <= 0.994105383;
cosLookup[1134] <= 0.994094983;
cosLookup[1135] <= 0.994084575;
cosLookup[1136] <= 0.994074157;
cosLookup[1137] <= 0.99406373;
cosLookup[1138] <= 0.994053293;
cosLookup[1139] <= 0.994042848;
cosLookup[1140] <= 0.994032394;
cosLookup[1141] <= 0.99402193;
cosLookup[1142] <= 0.994011457;
cosLookup[1143] <= 0.994000975;
cosLookup[1144] <= 0.993990484;
cosLookup[1145] <= 0.993979984;
cosLookup[1146] <= 0.993969475;
cosLookup[1147] <= 0.993958956;
cosLookup[1148] <= 0.993948429;
cosLookup[1149] <= 0.993937892;
cosLookup[1150] <= 0.993927346;
cosLookup[1151] <= 0.993916791;
cosLookup[1152] <= 0.993906227;
cosLookup[1153] <= 0.993895654;
cosLookup[1154] <= 0.993885071;
cosLookup[1155] <= 0.99387448;
cosLookup[1156] <= 0.993863879;
cosLookup[1157] <= 0.993853269;
cosLookup[1158] <= 0.99384265;
cosLookup[1159] <= 0.993832022;
cosLookup[1160] <= 0.993821385;
cosLookup[1161] <= 0.993810738;
cosLookup[1162] <= 0.993800083;
cosLookup[1163] <= 0.993789418;
cosLookup[1164] <= 0.993778745;
cosLookup[1165] <= 0.993768062;
cosLookup[1166] <= 0.99375737;
cosLookup[1167] <= 0.993746668;
cosLookup[1168] <= 0.993735958;
cosLookup[1169] <= 0.993725239;
cosLookup[1170] <= 0.99371451;
cosLookup[1171] <= 0.993703772;
cosLookup[1172] <= 0.993693025;
cosLookup[1173] <= 0.993682269;
cosLookup[1174] <= 0.993671504;
cosLookup[1175] <= 0.99366073;
cosLookup[1176] <= 0.993649947;
cosLookup[1177] <= 0.993639154;
cosLookup[1178] <= 0.993628352;
cosLookup[1179] <= 0.993617542;
cosLookup[1180] <= 0.993606722;
cosLookup[1181] <= 0.993595893;
cosLookup[1182] <= 0.993585054;
cosLookup[1183] <= 0.993574207;
cosLookup[1184] <= 0.993563351;
cosLookup[1185] <= 0.993552485;
cosLookup[1186] <= 0.99354161;
cosLookup[1187] <= 0.993530726;
cosLookup[1188] <= 0.993519833;
cosLookup[1189] <= 0.993508931;
cosLookup[1190] <= 0.99349802;
cosLookup[1191] <= 0.9934871;
cosLookup[1192] <= 0.99347617;
cosLookup[1193] <= 0.993465231;
cosLookup[1194] <= 0.993454284;
cosLookup[1195] <= 0.993443327;
cosLookup[1196] <= 0.993432361;
cosLookup[1197] <= 0.993421385;
cosLookup[1198] <= 0.993410401;
cosLookup[1199] <= 0.993399408;
cosLookup[1200] <= 0.993388405;
cosLookup[1201] <= 0.993377393;
cosLookup[1202] <= 0.993366372;
cosLookup[1203] <= 0.993355342;
cosLookup[1204] <= 0.993344303;
cosLookup[1205] <= 0.993333255;
cosLookup[1206] <= 0.993322198;
cosLookup[1207] <= 0.993311131;
cosLookup[1208] <= 0.993300055;
cosLookup[1209] <= 0.993288971;
cosLookup[1210] <= 0.993277877;
cosLookup[1211] <= 0.993266774;
cosLookup[1212] <= 0.993255662;
cosLookup[1213] <= 0.99324454;
cosLookup[1214] <= 0.99323341;
cosLookup[1215] <= 0.99322227;
cosLookup[1216] <= 0.993211121;
cosLookup[1217] <= 0.993199964;
cosLookup[1218] <= 0.993188797;
cosLookup[1219] <= 0.993177621;
cosLookup[1220] <= 0.993166435;
cosLookup[1221] <= 0.993155241;
cosLookup[1222] <= 0.993144038;
cosLookup[1223] <= 0.993132825;
cosLookup[1224] <= 0.993121603;
cosLookup[1225] <= 0.993110372;
cosLookup[1226] <= 0.993099132;
cosLookup[1227] <= 0.993087883;
cosLookup[1228] <= 0.993076625;
cosLookup[1229] <= 0.993065358;
cosLookup[1230] <= 0.993054081;
cosLookup[1231] <= 0.993042795;
cosLookup[1232] <= 0.993031501;
cosLookup[1233] <= 0.993020197;
cosLookup[1234] <= 0.993008884;
cosLookup[1235] <= 0.992997561;
cosLookup[1236] <= 0.99298623;
cosLookup[1237] <= 0.99297489;
cosLookup[1238] <= 0.99296354;
cosLookup[1239] <= 0.992952182;
cosLookup[1240] <= 0.992940814;
cosLookup[1241] <= 0.992929437;
cosLookup[1242] <= 0.992918051;
cosLookup[1243] <= 0.992906656;
cosLookup[1244] <= 0.992895251;
cosLookup[1245] <= 0.992883838;
cosLookup[1246] <= 0.992872415;
cosLookup[1247] <= 0.992860983;
cosLookup[1248] <= 0.992849543;
cosLookup[1249] <= 0.992838093;
cosLookup[1250] <= 0.992826634;
cosLookup[1251] <= 0.992815165;
cosLookup[1252] <= 0.992803688;
cosLookup[1253] <= 0.992792202;
cosLookup[1254] <= 0.992780706;
cosLookup[1255] <= 0.992769201;
cosLookup[1256] <= 0.992757687;
cosLookup[1257] <= 0.992746165;
cosLookup[1258] <= 0.992734632;
cosLookup[1259] <= 0.992723091;
cosLookup[1260] <= 0.992711541;
cosLookup[1261] <= 0.992699981;
cosLookup[1262] <= 0.992688413;
cosLookup[1263] <= 0.992676835;
cosLookup[1264] <= 0.992665248;
cosLookup[1265] <= 0.992653652;
cosLookup[1266] <= 0.992642047;
cosLookup[1267] <= 0.992630433;
cosLookup[1268] <= 0.99261881;
cosLookup[1269] <= 0.992607177;
cosLookup[1270] <= 0.992595535;
cosLookup[1271] <= 0.992583885;
cosLookup[1272] <= 0.992572225;
cosLookup[1273] <= 0.992560556;
cosLookup[1274] <= 0.992548878;
cosLookup[1275] <= 0.992537191;
cosLookup[1276] <= 0.992525494;
cosLookup[1277] <= 0.992513789;
cosLookup[1278] <= 0.992502074;
cosLookup[1279] <= 0.99249035;
cosLookup[1280] <= 0.992478618;
cosLookup[1281] <= 0.992466876;
cosLookup[1282] <= 0.992455125;
cosLookup[1283] <= 0.992443364;
cosLookup[1284] <= 0.992431595;
cosLookup[1285] <= 0.992419817;
cosLookup[1286] <= 0.992408029;
cosLookup[1287] <= 0.992396232;
cosLookup[1288] <= 0.992384426;
cosLookup[1289] <= 0.992372611;
cosLookup[1290] <= 0.992360787;
cosLookup[1291] <= 0.992348954;
cosLookup[1292] <= 0.992337112;
cosLookup[1293] <= 0.99232526;
cosLookup[1294] <= 0.9923134;
cosLookup[1295] <= 0.99230153;
cosLookup[1296] <= 0.992289651;
cosLookup[1297] <= 0.992277763;
cosLookup[1298] <= 0.992265866;
cosLookup[1299] <= 0.99225396;
cosLookup[1300] <= 0.992242045;
cosLookup[1301] <= 0.992230121;
cosLookup[1302] <= 0.992218187;
cosLookup[1303] <= 0.992206244;
cosLookup[1304] <= 0.992194293;
cosLookup[1305] <= 0.992182332;
cosLookup[1306] <= 0.992170362;
cosLookup[1307] <= 0.992158382;
cosLookup[1308] <= 0.992146394;
cosLookup[1309] <= 0.992134397;
cosLookup[1310] <= 0.99212239;
cosLookup[1311] <= 0.992110375;
cosLookup[1312] <= 0.99209835;
cosLookup[1313] <= 0.992086316;
cosLookup[1314] <= 0.992074273;
cosLookup[1315] <= 0.992062221;
cosLookup[1316] <= 0.99205016;
cosLookup[1317] <= 0.992038089;
cosLookup[1318] <= 0.99202601;
cosLookup[1319] <= 0.992013921;
cosLookup[1320] <= 0.992001824;
cosLookup[1321] <= 0.991989717;
cosLookup[1322] <= 0.991977601;
cosLookup[1323] <= 0.991965476;
cosLookup[1324] <= 0.991953342;
cosLookup[1325] <= 0.991941198;
cosLookup[1326] <= 0.991929046;
cosLookup[1327] <= 0.991916884;
cosLookup[1328] <= 0.991904714;
cosLookup[1329] <= 0.991892534;
cosLookup[1330] <= 0.991880345;
cosLookup[1331] <= 0.991868147;
cosLookup[1332] <= 0.99185594;
cosLookup[1333] <= 0.991843724;
cosLookup[1334] <= 0.991831498;
cosLookup[1335] <= 0.991819264;
cosLookup[1336] <= 0.99180702;
cosLookup[1337] <= 0.991794767;
cosLookup[1338] <= 0.991782505;
cosLookup[1339] <= 0.991770235;
cosLookup[1340] <= 0.991757954;
cosLookup[1341] <= 0.991745665;
cosLookup[1342] <= 0.991733367;
cosLookup[1343] <= 0.99172106;
cosLookup[1344] <= 0.991708743;
cosLookup[1345] <= 0.991696417;
cosLookup[1346] <= 0.991684083;
cosLookup[1347] <= 0.991671739;
cosLookup[1348] <= 0.991659386;
cosLookup[1349] <= 0.991647024;
cosLookup[1350] <= 0.991634652;
cosLookup[1351] <= 0.991622272;
cosLookup[1352] <= 0.991609882;
cosLookup[1353] <= 0.991597484;
cosLookup[1354] <= 0.991585076;
cosLookup[1355] <= 0.991572659;
cosLookup[1356] <= 0.991560233;
cosLookup[1357] <= 0.991547798;
cosLookup[1358] <= 0.991535354;
cosLookup[1359] <= 0.991522901;
cosLookup[1360] <= 0.991510438;
cosLookup[1361] <= 0.991497967;
cosLookup[1362] <= 0.991485486;
cosLookup[1363] <= 0.991472997;
cosLookup[1364] <= 0.991460498;
cosLookup[1365] <= 0.99144799;
cosLookup[1366] <= 0.991435473;
cosLookup[1367] <= 0.991422947;
cosLookup[1368] <= 0.991410411;
cosLookup[1369] <= 0.991397867;
cosLookup[1370] <= 0.991385313;
cosLookup[1371] <= 0.991372751;
cosLookup[1372] <= 0.991360179;
cosLookup[1373] <= 0.991347598;
cosLookup[1374] <= 0.991335008;
cosLookup[1375] <= 0.991322409;
cosLookup[1376] <= 0.991309801;
cosLookup[1377] <= 0.991297183;
cosLookup[1378] <= 0.991284557;
cosLookup[1379] <= 0.991271921;
cosLookup[1380] <= 0.991259277;
cosLookup[1381] <= 0.991246623;
cosLookup[1382] <= 0.99123396;
cosLookup[1383] <= 0.991221288;
cosLookup[1384] <= 0.991208607;
cosLookup[1385] <= 0.991195917;
cosLookup[1386] <= 0.991183217;
cosLookup[1387] <= 0.991170509;
cosLookup[1388] <= 0.991157791;
cosLookup[1389] <= 0.991145064;
cosLookup[1390] <= 0.991132329;
cosLookup[1391] <= 0.991119584;
cosLookup[1392] <= 0.99110683;
cosLookup[1393] <= 0.991094067;
cosLookup[1394] <= 0.991081294;
cosLookup[1395] <= 0.991068513;
cosLookup[1396] <= 0.991055723;
cosLookup[1397] <= 0.991042923;
cosLookup[1398] <= 0.991030114;
cosLookup[1399] <= 0.991017297;
cosLookup[1400] <= 0.99100447;
cosLookup[1401] <= 0.990991634;
cosLookup[1402] <= 0.990978789;
cosLookup[1403] <= 0.990965934;
cosLookup[1404] <= 0.990953071;
cosLookup[1405] <= 0.990940199;
cosLookup[1406] <= 0.990927317;
cosLookup[1407] <= 0.990914426;
cosLookup[1408] <= 0.990901526;
cosLookup[1409] <= 0.990888618;
cosLookup[1410] <= 0.9908757;
cosLookup[1411] <= 0.990862773;
cosLookup[1412] <= 0.990849836;
cosLookup[1413] <= 0.990836891;
cosLookup[1414] <= 0.990823937;
cosLookup[1415] <= 0.990810973;
cosLookup[1416] <= 0.990798;
cosLookup[1417] <= 0.990785019;
cosLookup[1418] <= 0.990772028;
cosLookup[1419] <= 0.990759028;
cosLookup[1420] <= 0.990746019;
cosLookup[1421] <= 0.990733;
cosLookup[1422] <= 0.990719973;
cosLookup[1423] <= 0.990706937;
cosLookup[1424] <= 0.990693891;
cosLookup[1425] <= 0.990680837;
cosLookup[1426] <= 0.990667773;
cosLookup[1427] <= 0.9906547;
cosLookup[1428] <= 0.990641618;
cosLookup[1429] <= 0.990628527;
cosLookup[1430] <= 0.990615427;
cosLookup[1431] <= 0.990602318;
cosLookup[1432] <= 0.990589199;
cosLookup[1433] <= 0.990576072;
cosLookup[1434] <= 0.990562935;
cosLookup[1435] <= 0.99054979;
cosLookup[1436] <= 0.990536635;
cosLookup[1437] <= 0.990523471;
cosLookup[1438] <= 0.990510298;
cosLookup[1439] <= 0.990497116;
cosLookup[1440] <= 0.990483925;
cosLookup[1441] <= 0.990470724;
cosLookup[1442] <= 0.990457515;
cosLookup[1443] <= 0.990444296;
cosLookup[1444] <= 0.990431069;
cosLookup[1445] <= 0.990417832;
cosLookup[1446] <= 0.990404586;
cosLookup[1447] <= 0.990391331;
cosLookup[1448] <= 0.990378067;
cosLookup[1449] <= 0.990364794;
cosLookup[1450] <= 0.990351512;
cosLookup[1451] <= 0.99033822;
cosLookup[1452] <= 0.99032492;
cosLookup[1453] <= 0.99031161;
cosLookup[1454] <= 0.990298291;
cosLookup[1455] <= 0.990284964;
cosLookup[1456] <= 0.990271627;
cosLookup[1457] <= 0.990258281;
cosLookup[1458] <= 0.990244926;
cosLookup[1459] <= 0.990231561;
cosLookup[1460] <= 0.990218188;
cosLookup[1461] <= 0.990204806;
cosLookup[1462] <= 0.990191414;
cosLookup[1463] <= 0.990178014;
cosLookup[1464] <= 0.990164604;
cosLookup[1465] <= 0.990151185;
cosLookup[1466] <= 0.990137757;
cosLookup[1467] <= 0.99012432;
cosLookup[1468] <= 0.990110874;
cosLookup[1469] <= 0.990097419;
cosLookup[1470] <= 0.990083955;
cosLookup[1471] <= 0.990070481;
cosLookup[1472] <= 0.990056999;
cosLookup[1473] <= 0.990043507;
cosLookup[1474] <= 0.990030006;
cosLookup[1475] <= 0.990016496;
cosLookup[1476] <= 0.990002977;
cosLookup[1477] <= 0.989989449;
cosLookup[1478] <= 0.989975912;
cosLookup[1479] <= 0.989962366;
cosLookup[1480] <= 0.989948811;
cosLookup[1481] <= 0.989935246;
cosLookup[1482] <= 0.989921673;
cosLookup[1483] <= 0.98990809;
cosLookup[1484] <= 0.989894498;
cosLookup[1485] <= 0.989880897;
cosLookup[1486] <= 0.989867288;
cosLookup[1487] <= 0.989853669;
cosLookup[1488] <= 0.98984004;
cosLookup[1489] <= 0.989826403;
cosLookup[1490] <= 0.989812757;
cosLookup[1491] <= 0.989799101;
cosLookup[1492] <= 0.989785437;
cosLookup[1493] <= 0.989771763;
cosLookup[1494] <= 0.98975808;
cosLookup[1495] <= 0.989744389;
cosLookup[1496] <= 0.989730688;
cosLookup[1497] <= 0.989716978;
cosLookup[1498] <= 0.989703259;
cosLookup[1499] <= 0.98968953;
cosLookup[1500] <= 0.989675793;
cosLookup[1501] <= 0.989662047;
cosLookup[1502] <= 0.989648291;
cosLookup[1503] <= 0.989634526;
cosLookup[1504] <= 0.989620753;
cosLookup[1505] <= 0.98960697;
cosLookup[1506] <= 0.989593178;
cosLookup[1507] <= 0.989579377;
cosLookup[1508] <= 0.989565567;
cosLookup[1509] <= 0.989551748;
cosLookup[1510] <= 0.989537919;
cosLookup[1511] <= 0.989524082;
cosLookup[1512] <= 0.989510235;
cosLookup[1513] <= 0.98949638;
cosLookup[1514] <= 0.989482515;
cosLookup[1515] <= 0.989468641;
cosLookup[1516] <= 0.989454759;
cosLookup[1517] <= 0.989440867;
cosLookup[1518] <= 0.989426965;
cosLookup[1519] <= 0.989413055;
cosLookup[1520] <= 0.989399136;
cosLookup[1521] <= 0.989385208;
cosLookup[1522] <= 0.98937127;
cosLookup[1523] <= 0.989357324;
cosLookup[1524] <= 0.989343368;
cosLookup[1525] <= 0.989329403;
cosLookup[1526] <= 0.98931543;
cosLookup[1527] <= 0.989301447;
cosLookup[1528] <= 0.989287455;
cosLookup[1529] <= 0.989273453;
cosLookup[1530] <= 0.989259443;
cosLookup[1531] <= 0.989245424;
cosLookup[1532] <= 0.989231396;
cosLookup[1533] <= 0.989217358;
cosLookup[1534] <= 0.989203311;
cosLookup[1535] <= 0.989189256;
cosLookup[1536] <= 0.989175191;
cosLookup[1537] <= 0.989161117;
cosLookup[1538] <= 0.989147034;
cosLookup[1539] <= 0.989132942;
cosLookup[1540] <= 0.989118841;
cosLookup[1541] <= 0.989104731;
cosLookup[1542] <= 0.989090611;
cosLookup[1543] <= 0.989076483;
cosLookup[1544] <= 0.989062345;
cosLookup[1545] <= 0.989048199;
cosLookup[1546] <= 0.989034043;
cosLookup[1547] <= 0.989019878;
cosLookup[1548] <= 0.989005704;
cosLookup[1549] <= 0.988991522;
cosLookup[1550] <= 0.988977329;
cosLookup[1551] <= 0.988963128;
cosLookup[1552] <= 0.988948918;
cosLookup[1553] <= 0.988934699;
cosLookup[1554] <= 0.98892047;
cosLookup[1555] <= 0.988906233;
cosLookup[1556] <= 0.988891986;
cosLookup[1557] <= 0.98887773;
cosLookup[1558] <= 0.988863466;
cosLookup[1559] <= 0.988849192;
cosLookup[1560] <= 0.988834909;
cosLookup[1561] <= 0.988820617;
cosLookup[1562] <= 0.988806316;
cosLookup[1563] <= 0.988792005;
cosLookup[1564] <= 0.988777686;
cosLookup[1565] <= 0.988763358;
cosLookup[1566] <= 0.98874902;
cosLookup[1567] <= 0.988734673;
cosLookup[1568] <= 0.988720318;
cosLookup[1569] <= 0.988705953;
cosLookup[1570] <= 0.988691579;
cosLookup[1571] <= 0.988677196;
cosLookup[1572] <= 0.988662804;
cosLookup[1573] <= 0.988648403;
cosLookup[1574] <= 0.988633993;
cosLookup[1575] <= 0.988619573;
cosLookup[1576] <= 0.988605145;
cosLookup[1577] <= 0.988590707;
cosLookup[1578] <= 0.988576261;
cosLookup[1579] <= 0.988561805;
cosLookup[1580] <= 0.98854734;
cosLookup[1581] <= 0.988532867;
cosLookup[1582] <= 0.988518384;
cosLookup[1583] <= 0.988503892;
cosLookup[1584] <= 0.98848939;
cosLookup[1585] <= 0.98847488;
cosLookup[1586] <= 0.988460361;
cosLookup[1587] <= 0.988445833;
cosLookup[1588] <= 0.988431295;
cosLookup[1589] <= 0.988416749;
cosLookup[1590] <= 0.988402193;
cosLookup[1591] <= 0.988387628;
cosLookup[1592] <= 0.988373055;
cosLookup[1593] <= 0.988358472;
cosLookup[1594] <= 0.98834388;
cosLookup[1595] <= 0.988329279;
cosLookup[1596] <= 0.988314668;
cosLookup[1597] <= 0.988300049;
cosLookup[1598] <= 0.988285421;
cosLookup[1599] <= 0.988270783;
cosLookup[1600] <= 0.988256137;
cosLookup[1601] <= 0.988241481;
cosLookup[1602] <= 0.988226817;
cosLookup[1603] <= 0.988212143;
cosLookup[1604] <= 0.98819746;
cosLookup[1605] <= 0.988182768;
cosLookup[1606] <= 0.988168067;
cosLookup[1607] <= 0.988153357;
cosLookup[1608] <= 0.988138638;
cosLookup[1609] <= 0.98812391;
cosLookup[1610] <= 0.988109173;
cosLookup[1611] <= 0.988094426;
cosLookup[1612] <= 0.988079671;
cosLookup[1613] <= 0.988064906;
cosLookup[1614] <= 0.988050132;
cosLookup[1615] <= 0.98803535;
cosLookup[1616] <= 0.988020558;
cosLookup[1617] <= 0.988005757;
cosLookup[1618] <= 0.987990947;
cosLookup[1619] <= 0.987976128;
cosLookup[1620] <= 0.9879613;
cosLookup[1621] <= 0.987946462;
cosLookup[1622] <= 0.987931616;
cosLookup[1623] <= 0.987916761;
cosLookup[1624] <= 0.987901896;
cosLookup[1625] <= 0.987887023;
cosLookup[1626] <= 0.98787214;
cosLookup[1627] <= 0.987857248;
cosLookup[1628] <= 0.987842347;
cosLookup[1629] <= 0.987827438;
cosLookup[1630] <= 0.987812519;
cosLookup[1631] <= 0.98779759;
cosLookup[1632] <= 0.987782653;
cosLookup[1633] <= 0.987767707;
cosLookup[1634] <= 0.987752752;
cosLookup[1635] <= 0.987737787;
cosLookup[1636] <= 0.987722814;
cosLookup[1637] <= 0.987707831;
cosLookup[1638] <= 0.98769284;
cosLookup[1639] <= 0.987677839;
cosLookup[1640] <= 0.987662829;
cosLookup[1641] <= 0.987647811;
cosLookup[1642] <= 0.987632783;
cosLookup[1643] <= 0.987617746;
cosLookup[1644] <= 0.987602699;
cosLookup[1645] <= 0.987587644;
cosLookup[1646] <= 0.98757258;
cosLookup[1647] <= 0.987557507;
cosLookup[1648] <= 0.987542424;
cosLookup[1649] <= 0.987527333;
cosLookup[1650] <= 0.987512232;
cosLookup[1651] <= 0.987497123;
cosLookup[1652] <= 0.987482004;
cosLookup[1653] <= 0.987466876;
cosLookup[1654] <= 0.987451739;
cosLookup[1655] <= 0.987436593;
cosLookup[1656] <= 0.987421438;
cosLookup[1657] <= 0.987406274;
cosLookup[1658] <= 0.987391101;
cosLookup[1659] <= 0.987375919;
cosLookup[1660] <= 0.987360727;
cosLookup[1661] <= 0.987345527;
cosLookup[1662] <= 0.987330317;
cosLookup[1663] <= 0.987315099;
cosLookup[1664] <= 0.987299871;
cosLookup[1665] <= 0.987284634;
cosLookup[1666] <= 0.987269389;
cosLookup[1667] <= 0.987254134;
cosLookup[1668] <= 0.98723887;
cosLookup[1669] <= 0.987223597;
cosLookup[1670] <= 0.987208315;
cosLookup[1671] <= 0.987193024;
cosLookup[1672] <= 0.987177723;
cosLookup[1673] <= 0.987162414;
cosLookup[1674] <= 0.987147096;
cosLookup[1675] <= 0.987131768;
cosLookup[1676] <= 0.987116432;
cosLookup[1677] <= 0.987101086;
cosLookup[1678] <= 0.987085731;
cosLookup[1679] <= 0.987070367;
cosLookup[1680] <= 0.987054995;
cosLookup[1681] <= 0.987039613;
cosLookup[1682] <= 0.987024222;
cosLookup[1683] <= 0.987008822;
cosLookup[1684] <= 0.986993412;
cosLookup[1685] <= 0.986977994;
cosLookup[1686] <= 0.986962567;
cosLookup[1687] <= 0.986947131;
cosLookup[1688] <= 0.986931685;
cosLookup[1689] <= 0.986916231;
cosLookup[1690] <= 0.986900767;
cosLookup[1691] <= 0.986885294;
cosLookup[1692] <= 0.986869813;
cosLookup[1693] <= 0.986854322;
cosLookup[1694] <= 0.986838822;
cosLookup[1695] <= 0.986823313;
cosLookup[1696] <= 0.986807795;
cosLookup[1697] <= 0.986792268;
cosLookup[1698] <= 0.986776732;
cosLookup[1699] <= 0.986761187;
cosLookup[1700] <= 0.986745632;
cosLookup[1701] <= 0.986730069;
cosLookup[1702] <= 0.986714496;
cosLookup[1703] <= 0.986698915;
cosLookup[1704] <= 0.986683324;
cosLookup[1705] <= 0.986667725;
cosLookup[1706] <= 0.986652116;
cosLookup[1707] <= 0.986636498;
cosLookup[1708] <= 0.986620871;
cosLookup[1709] <= 0.986605235;
cosLookup[1710] <= 0.98658959;
cosLookup[1711] <= 0.986573936;
cosLookup[1712] <= 0.986558273;
cosLookup[1713] <= 0.986542601;
cosLookup[1714] <= 0.98652692;
cosLookup[1715] <= 0.986511229;
cosLookup[1716] <= 0.98649553;
cosLookup[1717] <= 0.986479821;
cosLookup[1718] <= 0.986464104;
cosLookup[1719] <= 0.986448377;
cosLookup[1720] <= 0.986432642;
cosLookup[1721] <= 0.986416897;
cosLookup[1722] <= 0.986401143;
cosLookup[1723] <= 0.98638538;
cosLookup[1724] <= 0.986369608;
cosLookup[1725] <= 0.986353827;
cosLookup[1726] <= 0.986338037;
cosLookup[1727] <= 0.986322238;
cosLookup[1728] <= 0.98630643;
cosLookup[1729] <= 0.986290612;
cosLookup[1730] <= 0.986274786;
cosLookup[1731] <= 0.98625895;
cosLookup[1732] <= 0.986243106;
cosLookup[1733] <= 0.986227252;
cosLookup[1734] <= 0.98621139;
cosLookup[1735] <= 0.986195518;
cosLookup[1736] <= 0.986179637;
cosLookup[1737] <= 0.986163747;
cosLookup[1738] <= 0.986147849;
cosLookup[1739] <= 0.986131941;
cosLookup[1740] <= 0.986116024;
cosLookup[1741] <= 0.986100097;
cosLookup[1742] <= 0.986084162;
cosLookup[1743] <= 0.986068218;
cosLookup[1744] <= 0.986052265;
cosLookup[1745] <= 0.986036302;
cosLookup[1746] <= 0.986020331;
cosLookup[1747] <= 0.986004351;
cosLookup[1748] <= 0.985988361;
cosLookup[1749] <= 0.985972362;
cosLookup[1750] <= 0.985956355;
cosLookup[1751] <= 0.985940338;
cosLookup[1752] <= 0.985924312;
cosLookup[1753] <= 0.985908277;
cosLookup[1754] <= 0.985892233;
cosLookup[1755] <= 0.98587618;
cosLookup[1756] <= 0.985860118;
cosLookup[1757] <= 0.985844047;
cosLookup[1758] <= 0.985827967;
cosLookup[1759] <= 0.985811878;
cosLookup[1760] <= 0.985795779;
cosLookup[1761] <= 0.985779672;
cosLookup[1762] <= 0.985763556;
cosLookup[1763] <= 0.98574743;
cosLookup[1764] <= 0.985731296;
cosLookup[1765] <= 0.985715152;
cosLookup[1766] <= 0.985698999;
cosLookup[1767] <= 0.985682838;
cosLookup[1768] <= 0.985666667;
cosLookup[1769] <= 0.985650487;
cosLookup[1770] <= 0.985634298;
cosLookup[1771] <= 0.9856181;
cosLookup[1772] <= 0.985601893;
cosLookup[1773] <= 0.985585677;
cosLookup[1774] <= 0.985569452;
cosLookup[1775] <= 0.985553217;
cosLookup[1776] <= 0.985536974;
cosLookup[1777] <= 0.985520722;
cosLookup[1778] <= 0.98550446;
cosLookup[1779] <= 0.98548819;
cosLookup[1780] <= 0.98547191;
cosLookup[1781] <= 0.985455622;
cosLookup[1782] <= 0.985439324;
cosLookup[1783] <= 0.985423017;
cosLookup[1784] <= 0.985406702;
cosLookup[1785] <= 0.985390377;
cosLookup[1786] <= 0.985374043;
cosLookup[1787] <= 0.9853577;
cosLookup[1788] <= 0.985341348;
cosLookup[1789] <= 0.985324987;
cosLookup[1790] <= 0.985308617;
cosLookup[1791] <= 0.985292238;
cosLookup[1792] <= 0.985275849;
cosLookup[1793] <= 0.985259452;
cosLookup[1794] <= 0.985243046;
cosLookup[1795] <= 0.98522663;
cosLookup[1796] <= 0.985210206;
cosLookup[1797] <= 0.985193772;
cosLookup[1798] <= 0.98517733;
cosLookup[1799] <= 0.985160878;
cosLookup[1800] <= 0.985144418;
cosLookup[1801] <= 0.985127948;
cosLookup[1802] <= 0.985111469;
cosLookup[1803] <= 0.985094981;
cosLookup[1804] <= 0.985078484;
cosLookup[1805] <= 0.985061978;
cosLookup[1806] <= 0.985045463;
cosLookup[1807] <= 0.985028939;
cosLookup[1808] <= 0.985012406;
cosLookup[1809] <= 0.984995864;
cosLookup[1810] <= 0.984979313;
cosLookup[1811] <= 0.984962752;
cosLookup[1812] <= 0.984946183;
cosLookup[1813] <= 0.984929605;
cosLookup[1814] <= 0.984913017;
cosLookup[1815] <= 0.984896421;
cosLookup[1816] <= 0.984879815;
cosLookup[1817] <= 0.9848632;
cosLookup[1818] <= 0.984846577;
cosLookup[1819] <= 0.984829944;
cosLookup[1820] <= 0.984813302;
cosLookup[1821] <= 0.984796651;
cosLookup[1822] <= 0.984779992;
cosLookup[1823] <= 0.984763323;
cosLookup[1824] <= 0.984746645;
cosLookup[1825] <= 0.984729958;
cosLookup[1826] <= 0.984713261;
cosLookup[1827] <= 0.984696556;
cosLookup[1828] <= 0.984679842;
cosLookup[1829] <= 0.984663119;
cosLookup[1830] <= 0.984646387;
cosLookup[1831] <= 0.984629645;
cosLookup[1832] <= 0.984612895;
cosLookup[1833] <= 0.984596135;
cosLookup[1834] <= 0.984579367;
cosLookup[1835] <= 0.984562589;
cosLookup[1836] <= 0.984545803;
cosLookup[1837] <= 0.984529007;
cosLookup[1838] <= 0.984512202;
cosLookup[1839] <= 0.984495388;
cosLookup[1840] <= 0.984478566;
cosLookup[1841] <= 0.984461734;
cosLookup[1842] <= 0.984444893;
cosLookup[1843] <= 0.984428043;
cosLookup[1844] <= 0.984411184;
cosLookup[1845] <= 0.984394316;
cosLookup[1846] <= 0.984377439;
cosLookup[1847] <= 0.984360553;
cosLookup[1848] <= 0.984343657;
cosLookup[1849] <= 0.984326753;
cosLookup[1850] <= 0.98430984;
cosLookup[1851] <= 0.984292917;
cosLookup[1852] <= 0.984275986;
cosLookup[1853] <= 0.984259045;
cosLookup[1854] <= 0.984242096;
cosLookup[1855] <= 0.984225137;
cosLookup[1856] <= 0.98420817;
cosLookup[1857] <= 0.984191193;
cosLookup[1858] <= 0.984174207;
cosLookup[1859] <= 0.984157213;
cosLookup[1860] <= 0.984140209;
cosLookup[1861] <= 0.984123196;
cosLookup[1862] <= 0.984106174;
cosLookup[1863] <= 0.984089143;
cosLookup[1864] <= 0.984072103;
cosLookup[1865] <= 0.984055054;
cosLookup[1866] <= 0.984037996;
cosLookup[1867] <= 0.984020929;
cosLookup[1868] <= 0.984003853;
cosLookup[1869] <= 0.983986768;
cosLookup[1870] <= 0.983969673;
cosLookup[1871] <= 0.98395257;
cosLookup[1872] <= 0.983935458;
cosLookup[1873] <= 0.983918336;
cosLookup[1874] <= 0.983901206;
cosLookup[1875] <= 0.983884066;
cosLookup[1876] <= 0.983866918;
cosLookup[1877] <= 0.98384976;
cosLookup[1878] <= 0.983832594;
cosLookup[1879] <= 0.983815418;
cosLookup[1880] <= 0.983798233;
cosLookup[1881] <= 0.98378104;
cosLookup[1882] <= 0.983763837;
cosLookup[1883] <= 0.983746625;
cosLookup[1884] <= 0.983729404;
cosLookup[1885] <= 0.983712174;
cosLookup[1886] <= 0.983694935;
cosLookup[1887] <= 0.983677687;
cosLookup[1888] <= 0.98366043;
cosLookup[1889] <= 0.983643164;
cosLookup[1890] <= 0.983625889;
cosLookup[1891] <= 0.983608605;
cosLookup[1892] <= 0.983591312;
cosLookup[1893] <= 0.983574009;
cosLookup[1894] <= 0.983556698;
cosLookup[1895] <= 0.983539378;
cosLookup[1896] <= 0.983522048;
cosLookup[1897] <= 0.98350471;
cosLookup[1898] <= 0.983487362;
cosLookup[1899] <= 0.983470006;
cosLookup[1900] <= 0.98345264;
cosLookup[1901] <= 0.983435266;
cosLookup[1902] <= 0.983417882;
cosLookup[1903] <= 0.983400489;
cosLookup[1904] <= 0.983383088;
cosLookup[1905] <= 0.983365677;
cosLookup[1906] <= 0.983348257;
cosLookup[1907] <= 0.983330828;
cosLookup[1908] <= 0.98331339;
cosLookup[1909] <= 0.983295943;
cosLookup[1910] <= 0.983278487;
cosLookup[1911] <= 0.983261022;
cosLookup[1912] <= 0.983243548;
cosLookup[1913] <= 0.983226065;
cosLookup[1914] <= 0.983208573;
cosLookup[1915] <= 0.983191072;
cosLookup[1916] <= 0.983173562;
cosLookup[1917] <= 0.983156043;
cosLookup[1918] <= 0.983138514;
cosLookup[1919] <= 0.983120977;
cosLookup[1920] <= 0.983103431;
cosLookup[1921] <= 0.983085875;
cosLookup[1922] <= 0.983068311;
cosLookup[1923] <= 0.983050738;
cosLookup[1924] <= 0.983033155;
cosLookup[1925] <= 0.983015563;
cosLookup[1926] <= 0.982997963;
cosLookup[1927] <= 0.982980353;
cosLookup[1928] <= 0.982962735;
cosLookup[1929] <= 0.982945107;
cosLookup[1930] <= 0.98292747;
cosLookup[1931] <= 0.982909825;
cosLookup[1932] <= 0.98289217;
cosLookup[1933] <= 0.982874506;
cosLookup[1934] <= 0.982856833;
cosLookup[1935] <= 0.982839151;
cosLookup[1936] <= 0.98282146;
cosLookup[1937] <= 0.98280376;
cosLookup[1938] <= 0.982786051;
cosLookup[1939] <= 0.982768333;
cosLookup[1940] <= 0.982750606;
cosLookup[1941] <= 0.98273287;
cosLookup[1942] <= 0.982715125;
cosLookup[1943] <= 0.982697371;
cosLookup[1944] <= 0.982679608;
cosLookup[1945] <= 0.982661835;
cosLookup[1946] <= 0.982644054;
cosLookup[1947] <= 0.982626264;
cosLookup[1948] <= 0.982608465;
cosLookup[1949] <= 0.982590656;
cosLookup[1950] <= 0.982572839;
cosLookup[1951] <= 0.982555012;
cosLookup[1952] <= 0.982537177;
cosLookup[1953] <= 0.982519332;
cosLookup[1954] <= 0.982501479;
cosLookup[1955] <= 0.982483616;
cosLookup[1956] <= 0.982465745;
cosLookup[1957] <= 0.982447864;
cosLookup[1958] <= 0.982429974;
cosLookup[1959] <= 0.982412076;
cosLookup[1960] <= 0.982394168;
cosLookup[1961] <= 0.982376251;
cosLookup[1962] <= 0.982358326;
cosLookup[1963] <= 0.982340391;
cosLookup[1964] <= 0.982322447;
cosLookup[1965] <= 0.982304494;
cosLookup[1966] <= 0.982286532;
cosLookup[1967] <= 0.982268561;
cosLookup[1968] <= 0.982250581;
cosLookup[1969] <= 0.982232592;
cosLookup[1970] <= 0.982214594;
cosLookup[1971] <= 0.982196587;
cosLookup[1972] <= 0.982178571;
cosLookup[1973] <= 0.982160546;
cosLookup[1974] <= 0.982142512;
cosLookup[1975] <= 0.982124469;
cosLookup[1976] <= 0.982106416;
cosLookup[1977] <= 0.982088355;
cosLookup[1978] <= 0.982070285;
cosLookup[1979] <= 0.982052206;
cosLookup[1980] <= 0.982034117;
cosLookup[1981] <= 0.98201602;
cosLookup[1982] <= 0.981997914;
cosLookup[1983] <= 0.981979798;
cosLookup[1984] <= 0.981961674;
cosLookup[1985] <= 0.98194354;
cosLookup[1986] <= 0.981925398;
cosLookup[1987] <= 0.981907246;
cosLookup[1988] <= 0.981889086;
cosLookup[1989] <= 0.981870916;
cosLookup[1990] <= 0.981852738;
cosLookup[1991] <= 0.98183455;
cosLookup[1992] <= 0.981816354;
cosLookup[1993] <= 0.981798148;
cosLookup[1994] <= 0.981779933;
cosLookup[1995] <= 0.98176171;
cosLookup[1996] <= 0.981743477;
cosLookup[1997] <= 0.981725235;
cosLookup[1998] <= 0.981706984;
cosLookup[1999] <= 0.981688724;
cosLookup[2000] <= 0.981670456;
cosLookup[2001] <= 0.981652178;
cosLookup[2002] <= 0.981633891;
cosLookup[2003] <= 0.981615595;
cosLookup[2004] <= 0.98159729;
cosLookup[2005] <= 0.981578976;
cosLookup[2006] <= 0.981560653;
cosLookup[2007] <= 0.981542321;
cosLookup[2008] <= 0.98152398;
cosLookup[2009] <= 0.98150563;
cosLookup[2010] <= 0.981487271;
cosLookup[2011] <= 0.981468903;
cosLookup[2012] <= 0.981450526;
cosLookup[2013] <= 0.98143214;
cosLookup[2014] <= 0.981413745;
cosLookup[2015] <= 0.98139534;
cosLookup[2016] <= 0.981376927;
cosLookup[2017] <= 0.981358505;
cosLookup[2018] <= 0.981340074;
cosLookup[2019] <= 0.981321633;
cosLookup[2020] <= 0.981303184;
cosLookup[2021] <= 0.981284726;
cosLookup[2022] <= 0.981266258;
cosLookup[2023] <= 0.981247782;
cosLookup[2024] <= 0.981229297;
cosLookup[2025] <= 0.981210802;
cosLookup[2026] <= 0.981192299;
cosLookup[2027] <= 0.981173787;
cosLookup[2028] <= 0.981155265;
cosLookup[2029] <= 0.981136735;
cosLookup[2030] <= 0.981118195;
cosLookup[2031] <= 0.981099647;
cosLookup[2032] <= 0.981081089;
cosLookup[2033] <= 0.981062523;
cosLookup[2034] <= 0.981043947;
cosLookup[2035] <= 0.981025362;
cosLookup[2036] <= 0.981006769;
cosLookup[2037] <= 0.980988166;
cosLookup[2038] <= 0.980969555;
cosLookup[2039] <= 0.980950934;
cosLookup[2040] <= 0.980932304;
cosLookup[2041] <= 0.980913666;
cosLookup[2042] <= 0.980895018;
cosLookup[2043] <= 0.980876361;
cosLookup[2044] <= 0.980857695;
cosLookup[2045] <= 0.980839021;
cosLookup[2046] <= 0.980820337;
cosLookup[2047] <= 0.980801644;
cosLookup[2048] <= 0.980782942;
cosLookup[2049] <= 0.980764231;
cosLookup[2050] <= 0.980745512;
cosLookup[2051] <= 0.980726783;
cosLookup[2052] <= 0.980708045;
cosLookup[2053] <= 0.980689298;
cosLookup[2054] <= 0.980670542;
cosLookup[2055] <= 0.980651777;
cosLookup[2056] <= 0.980633003;
cosLookup[2057] <= 0.98061422;
cosLookup[2058] <= 0.980595428;
cosLookup[2059] <= 0.980576627;
cosLookup[2060] <= 0.980557817;
cosLookup[2061] <= 0.980538998;
cosLookup[2062] <= 0.98052017;
cosLookup[2063] <= 0.980501333;
cosLookup[2064] <= 0.980482487;
cosLookup[2065] <= 0.980463632;
cosLookup[2066] <= 0.980444768;
cosLookup[2067] <= 0.980425895;
cosLookup[2068] <= 0.980407013;
cosLookup[2069] <= 0.980388122;
cosLookup[2070] <= 0.980369222;
cosLookup[2071] <= 0.980350312;
cosLookup[2072] <= 0.980331394;
cosLookup[2073] <= 0.980312467;
cosLookup[2074] <= 0.980293531;
cosLookup[2075] <= 0.980274586;
cosLookup[2076] <= 0.980255632;
cosLookup[2077] <= 0.980236668;
cosLookup[2078] <= 0.980217696;
cosLookup[2079] <= 0.980198715;
cosLookup[2080] <= 0.980179725;
cosLookup[2081] <= 0.980160725;
cosLookup[2082] <= 0.980141717;
cosLookup[2083] <= 0.9801227;
cosLookup[2084] <= 0.980103674;
cosLookup[2085] <= 0.980084638;
cosLookup[2086] <= 0.980065594;
cosLookup[2087] <= 0.980046541;
cosLookup[2088] <= 0.980027478;
cosLookup[2089] <= 0.980008407;
cosLookup[2090] <= 0.979989327;
cosLookup[2091] <= 0.979970237;
cosLookup[2092] <= 0.979951139;
cosLookup[2093] <= 0.979932032;
cosLookup[2094] <= 0.979912915;
cosLookup[2095] <= 0.97989379;
cosLookup[2096] <= 0.979874655;
cosLookup[2097] <= 0.979855512;
cosLookup[2098] <= 0.97983636;
cosLookup[2099] <= 0.979817198;
cosLookup[2100] <= 0.979798028;
cosLookup[2101] <= 0.979778848;
cosLookup[2102] <= 0.97975966;
cosLookup[2103] <= 0.979740462;
cosLookup[2104] <= 0.979721256;
cosLookup[2105] <= 0.97970204;
cosLookup[2106] <= 0.979682816;
cosLookup[2107] <= 0.979663583;
cosLookup[2108] <= 0.97964434;
cosLookup[2109] <= 0.979625089;
cosLookup[2110] <= 0.979605828;
cosLookup[2111] <= 0.979586559;
cosLookup[2112] <= 0.97956728;
cosLookup[2113] <= 0.979547993;
cosLookup[2114] <= 0.979528696;
cosLookup[2115] <= 0.979509391;
cosLookup[2116] <= 0.979490076;
cosLookup[2117] <= 0.979470752;
cosLookup[2118] <= 0.97945142;
cosLookup[2119] <= 0.979432078;
cosLookup[2120] <= 0.979412728;
cosLookup[2121] <= 0.979393368;
cosLookup[2122] <= 0.979374;
cosLookup[2123] <= 0.979354622;
cosLookup[2124] <= 0.979335236;
cosLookup[2125] <= 0.97931584;
cosLookup[2126] <= 0.979296436;
cosLookup[2127] <= 0.979277022;
cosLookup[2128] <= 0.979257599;
cosLookup[2129] <= 0.979238168;
cosLookup[2130] <= 0.979218727;
cosLookup[2131] <= 0.979199278;
cosLookup[2132] <= 0.979179819;
cosLookup[2133] <= 0.979160352;
cosLookup[2134] <= 0.979140875;
cosLookup[2135] <= 0.97912139;
cosLookup[2136] <= 0.979101895;
cosLookup[2137] <= 0.979082391;
cosLookup[2138] <= 0.979062879;
cosLookup[2139] <= 0.979043357;
cosLookup[2140] <= 0.979023827;
cosLookup[2141] <= 0.979004287;
cosLookup[2142] <= 0.978984738;
cosLookup[2143] <= 0.978965181;
cosLookup[2144] <= 0.978945614;
cosLookup[2145] <= 0.978926039;
cosLookup[2146] <= 0.978906454;
cosLookup[2147] <= 0.978886861;
cosLookup[2148] <= 0.978867258;
cosLookup[2149] <= 0.978847646;
cosLookup[2150] <= 0.978828026;
cosLookup[2151] <= 0.978808396;
cosLookup[2152] <= 0.978788758;
cosLookup[2153] <= 0.97876911;
cosLookup[2154] <= 0.978749454;
cosLookup[2155] <= 0.978729788;
cosLookup[2156] <= 0.978710114;
cosLookup[2157] <= 0.97869043;
cosLookup[2158] <= 0.978670737;
cosLookup[2159] <= 0.978651036;
cosLookup[2160] <= 0.978631325;
cosLookup[2161] <= 0.978611606;
cosLookup[2162] <= 0.978591877;
cosLookup[2163] <= 0.97857214;
cosLookup[2164] <= 0.978552393;
cosLookup[2165] <= 0.978532638;
cosLookup[2166] <= 0.978512873;
cosLookup[2167] <= 0.9784931;
cosLookup[2168] <= 0.978473317;
cosLookup[2169] <= 0.978453526;
cosLookup[2170] <= 0.978433725;
cosLookup[2171] <= 0.978413916;
cosLookup[2172] <= 0.978394097;
cosLookup[2173] <= 0.97837427;
cosLookup[2174] <= 0.978354433;
cosLookup[2175] <= 0.978334588;
cosLookup[2176] <= 0.978314733;
cosLookup[2177] <= 0.97829487;
cosLookup[2178] <= 0.978274997;
cosLookup[2179] <= 0.978255116;
cosLookup[2180] <= 0.978235225;
cosLookup[2181] <= 0.978215326;
cosLookup[2182] <= 0.978195418;
cosLookup[2183] <= 0.9781755;
cosLookup[2184] <= 0.978155574;
cosLookup[2185] <= 0.978135638;
cosLookup[2186] <= 0.978115694;
cosLookup[2187] <= 0.978095741;
cosLookup[2188] <= 0.978075778;
cosLookup[2189] <= 0.978055807;
cosLookup[2190] <= 0.978035827;
cosLookup[2191] <= 0.978015837;
cosLookup[2192] <= 0.977995839;
cosLookup[2193] <= 0.977975832;
cosLookup[2194] <= 0.977955815;
cosLookup[2195] <= 0.97793579;
cosLookup[2196] <= 0.977915756;
cosLookup[2197] <= 0.977895712;
cosLookup[2198] <= 0.97787566;
cosLookup[2199] <= 0.977855599;
cosLookup[2200] <= 0.977835528;
cosLookup[2201] <= 0.977815449;
cosLookup[2202] <= 0.977795361;
cosLookup[2203] <= 0.977775264;
cosLookup[2204] <= 0.977755158;
cosLookup[2205] <= 0.977735042;
cosLookup[2206] <= 0.977714918;
cosLookup[2207] <= 0.977694785;
cosLookup[2208] <= 0.977674643;
cosLookup[2209] <= 0.977654492;
cosLookup[2210] <= 0.977634332;
cosLookup[2211] <= 0.977614162;
cosLookup[2212] <= 0.977593984;
cosLookup[2213] <= 0.977573797;
cosLookup[2214] <= 0.977553601;
cosLookup[2215] <= 0.977533396;
cosLookup[2216] <= 0.977513182;
cosLookup[2217] <= 0.977492959;
cosLookup[2218] <= 0.977472727;
cosLookup[2219] <= 0.977452486;
cosLookup[2220] <= 0.977432236;
cosLookup[2221] <= 0.977411977;
cosLookup[2222] <= 0.977391709;
cosLookup[2223] <= 0.977371432;
cosLookup[2224] <= 0.977351146;
cosLookup[2225] <= 0.977330851;
cosLookup[2226] <= 0.977310547;
cosLookup[2227] <= 0.977290234;
cosLookup[2228] <= 0.977269912;
cosLookup[2229] <= 0.977249581;
cosLookup[2230] <= 0.977229242;
cosLookup[2231] <= 0.977208893;
cosLookup[2232] <= 0.977188535;
cosLookup[2233] <= 0.977168168;
cosLookup[2234] <= 0.977147792;
cosLookup[2235] <= 0.977127408;
cosLookup[2236] <= 0.977107014;
cosLookup[2237] <= 0.977086611;
cosLookup[2238] <= 0.977066199;
cosLookup[2239] <= 0.977045779;
cosLookup[2240] <= 0.977025349;
cosLookup[2241] <= 0.97700491;
cosLookup[2242] <= 0.976984463;
cosLookup[2243] <= 0.976964006;
cosLookup[2244] <= 0.97694354;
cosLookup[2245] <= 0.976923066;
cosLookup[2246] <= 0.976902582;
cosLookup[2247] <= 0.97688209;
cosLookup[2248] <= 0.976861588;
cosLookup[2249] <= 0.976841078;
cosLookup[2250] <= 0.976820558;
cosLookup[2251] <= 0.97680003;
cosLookup[2252] <= 0.976779492;
cosLookup[2253] <= 0.976758946;
cosLookup[2254] <= 0.97673839;
cosLookup[2255] <= 0.976717826;
cosLookup[2256] <= 0.976697253;
cosLookup[2257] <= 0.97667667;
cosLookup[2258] <= 0.976656079;
cosLookup[2259] <= 0.976635479;
cosLookup[2260] <= 0.976614869;
cosLookup[2261] <= 0.976594251;
cosLookup[2262] <= 0.976573624;
cosLookup[2263] <= 0.976552988;
cosLookup[2264] <= 0.976532343;
cosLookup[2265] <= 0.976511688;
cosLookup[2266] <= 0.976491025;
cosLookup[2267] <= 0.976470353;
cosLookup[2268] <= 0.976449672;
cosLookup[2269] <= 0.976428982;
cosLookup[2270] <= 0.976408283;
cosLookup[2271] <= 0.976387575;
cosLookup[2272] <= 0.976366858;
cosLookup[2273] <= 0.976346132;
cosLookup[2274] <= 0.976325397;
cosLookup[2275] <= 0.976304653;
cosLookup[2276] <= 0.9762839;
cosLookup[2277] <= 0.976263138;
cosLookup[2278] <= 0.976242367;
cosLookup[2279] <= 0.976221588;
cosLookup[2280] <= 0.976200799;
cosLookup[2281] <= 0.976180001;
cosLookup[2282] <= 0.976159194;
cosLookup[2283] <= 0.976138379;
cosLookup[2284] <= 0.976117554;
cosLookup[2285] <= 0.97609672;
cosLookup[2286] <= 0.976075878;
cosLookup[2287] <= 0.976055026;
cosLookup[2288] <= 0.976034165;
cosLookup[2289] <= 0.976013296;
cosLookup[2290] <= 0.975992417;
cosLookup[2291] <= 0.97597153;
cosLookup[2292] <= 0.975950633;
cosLookup[2293] <= 0.975929728;
cosLookup[2294] <= 0.975908813;
cosLookup[2295] <= 0.97588789;
cosLookup[2296] <= 0.975866958;
cosLookup[2297] <= 0.975846016;
cosLookup[2298] <= 0.975825066;
cosLookup[2299] <= 0.975804107;
cosLookup[2300] <= 0.975783138;
cosLookup[2301] <= 0.975762161;
cosLookup[2302] <= 0.975741175;
cosLookup[2303] <= 0.97572018;
cosLookup[2304] <= 0.975699176;
cosLookup[2305] <= 0.975678163;
cosLookup[2306] <= 0.975657141;
cosLookup[2307] <= 0.97563611;
cosLookup[2308] <= 0.97561507;
cosLookup[2309] <= 0.975594021;
cosLookup[2310] <= 0.975572963;
cosLookup[2311] <= 0.975551896;
cosLookup[2312] <= 0.97553082;
cosLookup[2313] <= 0.975509735;
cosLookup[2314] <= 0.975488641;
cosLookup[2315] <= 0.975467538;
cosLookup[2316] <= 0.975446427;
cosLookup[2317] <= 0.975425306;
cosLookup[2318] <= 0.975404176;
cosLookup[2319] <= 0.975383038;
cosLookup[2320] <= 0.97536189;
cosLookup[2321] <= 0.975340733;
cosLookup[2322] <= 0.975319568;
cosLookup[2323] <= 0.975298393;
cosLookup[2324] <= 0.97527721;
cosLookup[2325] <= 0.975256017;
cosLookup[2326] <= 0.975234816;
cosLookup[2327] <= 0.975213606;
cosLookup[2328] <= 0.975192386;
cosLookup[2329] <= 0.975171158;
cosLookup[2330] <= 0.975149921;
cosLookup[2331] <= 0.975128675;
cosLookup[2332] <= 0.975107419;
cosLookup[2333] <= 0.975086155;
cosLookup[2334] <= 0.975064882;
cosLookup[2335] <= 0.9750436;
cosLookup[2336] <= 0.975022309;
cosLookup[2337] <= 0.975001009;
cosLookup[2338] <= 0.9749797;
cosLookup[2339] <= 0.974958382;
cosLookup[2340] <= 0.974937055;
cosLookup[2341] <= 0.974915719;
cosLookup[2342] <= 0.974894374;
cosLookup[2343] <= 0.974873021;
cosLookup[2344] <= 0.974851658;
cosLookup[2345] <= 0.974830286;
cosLookup[2346] <= 0.974808905;
cosLookup[2347] <= 0.974787516;
cosLookup[2348] <= 0.974766117;
cosLookup[2349] <= 0.97474471;
cosLookup[2350] <= 0.974723293;
cosLookup[2351] <= 0.974701868;
cosLookup[2352] <= 0.974680433;
cosLookup[2353] <= 0.97465899;
cosLookup[2354] <= 0.974637537;
cosLookup[2355] <= 0.974616076;
cosLookup[2356] <= 0.974594606;
cosLookup[2357] <= 0.974573127;
cosLookup[2358] <= 0.974551638;
cosLookup[2359] <= 0.974530141;
cosLookup[2360] <= 0.974508635;
cosLookup[2361] <= 0.97448712;
cosLookup[2362] <= 0.974465596;
cosLookup[2363] <= 0.974444063;
cosLookup[2364] <= 0.974422521;
cosLookup[2365] <= 0.97440097;
cosLookup[2366] <= 0.97437941;
cosLookup[2367] <= 0.974357841;
cosLookup[2368] <= 0.974336264;
cosLookup[2369] <= 0.974314677;
cosLookup[2370] <= 0.974293081;
cosLookup[2371] <= 0.974271476;
cosLookup[2372] <= 0.974249863;
cosLookup[2373] <= 0.97422824;
cosLookup[2374] <= 0.974206609;
cosLookup[2375] <= 0.974184968;
cosLookup[2376] <= 0.974163319;
cosLookup[2377] <= 0.97414166;
cosLookup[2378] <= 0.974119993;
cosLookup[2379] <= 0.974098317;
cosLookup[2380] <= 0.974076632;
cosLookup[2381] <= 0.974054937;
cosLookup[2382] <= 0.974033234;
cosLookup[2383] <= 0.974011522;
cosLookup[2384] <= 0.973989801;
cosLookup[2385] <= 0.973968071;
cosLookup[2386] <= 0.973946332;
cosLookup[2387] <= 0.973924584;
cosLookup[2388] <= 0.973902827;
cosLookup[2389] <= 0.973881061;
cosLookup[2390] <= 0.973859287;
cosLookup[2391] <= 0.973837503;
cosLookup[2392] <= 0.97381571;
cosLookup[2393] <= 0.973793908;
cosLookup[2394] <= 0.973772098;
cosLookup[2395] <= 0.973750278;
cosLookup[2396] <= 0.97372845;
cosLookup[2397] <= 0.973706612;
cosLookup[2398] <= 0.973684766;
cosLookup[2399] <= 0.973662911;
cosLookup[2400] <= 0.973641046;
cosLookup[2401] <= 0.973619173;
cosLookup[2402] <= 0.973597291;
cosLookup[2403] <= 0.9735754;
cosLookup[2404] <= 0.9735535;
cosLookup[2405] <= 0.973531591;
cosLookup[2406] <= 0.973509673;
cosLookup[2407] <= 0.973487746;
cosLookup[2408] <= 0.97346581;
cosLookup[2409] <= 0.973443865;
cosLookup[2410] <= 0.973421911;
cosLookup[2411] <= 0.973399948;
cosLookup[2412] <= 0.973377977;
cosLookup[2413] <= 0.973355996;
cosLookup[2414] <= 0.973334006;
cosLookup[2415] <= 0.973312008;
cosLookup[2416] <= 0.97329;
cosLookup[2417] <= 0.973267984;
cosLookup[2418] <= 0.973245958;
cosLookup[2419] <= 0.973223924;
cosLookup[2420] <= 0.973201881;
cosLookup[2421] <= 0.973179829;
cosLookup[2422] <= 0.973157767;
cosLookup[2423] <= 0.973135697;
cosLookup[2424] <= 0.973113618;
cosLookup[2425] <= 0.97309153;
cosLookup[2426] <= 0.973069433;
cosLookup[2427] <= 0.973047327;
cosLookup[2428] <= 0.973025212;
cosLookup[2429] <= 0.973003089;
cosLookup[2430] <= 0.972980956;
cosLookup[2431] <= 0.972958814;
cosLookup[2432] <= 0.972936664;
cosLookup[2433] <= 0.972914504;
cosLookup[2434] <= 0.972892336;
cosLookup[2435] <= 0.972870158;
cosLookup[2436] <= 0.972847972;
cosLookup[2437] <= 0.972825776;
cosLookup[2438] <= 0.972803572;
cosLookup[2439] <= 0.972781359;
cosLookup[2440] <= 0.972759137;
cosLookup[2441] <= 0.972736906;
cosLookup[2442] <= 0.972714665;
cosLookup[2443] <= 0.972692416;
cosLookup[2444] <= 0.972670159;
cosLookup[2445] <= 0.972647892;
cosLookup[2446] <= 0.972625616;
cosLookup[2447] <= 0.972603331;
cosLookup[2448] <= 0.972581037;
cosLookup[2449] <= 0.972558735;
cosLookup[2450] <= 0.972536423;
cosLookup[2451] <= 0.972514103;
cosLookup[2452] <= 0.972491773;
cosLookup[2453] <= 0.972469435;
cosLookup[2454] <= 0.972447087;
cosLookup[2455] <= 0.972424731;
cosLookup[2456] <= 0.972402366;
cosLookup[2457] <= 0.972379992;
cosLookup[2458] <= 0.972357609;
cosLookup[2459] <= 0.972335217;
cosLookup[2460] <= 0.972312816;
cosLookup[2461] <= 0.972290406;
cosLookup[2462] <= 0.972267987;
cosLookup[2463] <= 0.972245559;
cosLookup[2464] <= 0.972223122;
cosLookup[2465] <= 0.972200677;
cosLookup[2466] <= 0.972178222;
cosLookup[2467] <= 0.972155758;
cosLookup[2468] <= 0.972133286;
cosLookup[2469] <= 0.972110804;
cosLookup[2470] <= 0.972088314;
cosLookup[2471] <= 0.972065815;
cosLookup[2472] <= 0.972043307;
cosLookup[2473] <= 0.972020789;
cosLookup[2474] <= 0.971998263;
cosLookup[2475] <= 0.971975728;
cosLookup[2476] <= 0.971953184;
cosLookup[2477] <= 0.971930631;
cosLookup[2478] <= 0.97190807;
cosLookup[2479] <= 0.971885499;
cosLookup[2480] <= 0.971862919;
cosLookup[2481] <= 0.97184033;
cosLookup[2482] <= 0.971817733;
cosLookup[2483] <= 0.971795126;
cosLookup[2484] <= 0.971772511;
cosLookup[2485] <= 0.971749887;
cosLookup[2486] <= 0.971727253;
cosLookup[2487] <= 0.971704611;
cosLookup[2488] <= 0.97168196;
cosLookup[2489] <= 0.9716593;
cosLookup[2490] <= 0.971636631;
cosLookup[2491] <= 0.971613953;
cosLookup[2492] <= 0.971591266;
cosLookup[2493] <= 0.97156857;
cosLookup[2494] <= 0.971545865;
cosLookup[2495] <= 0.971523151;
cosLookup[2496] <= 0.971500429;
cosLookup[2497] <= 0.971477697;
cosLookup[2498] <= 0.971454957;
cosLookup[2499] <= 0.971432207;
cosLookup[2500] <= 0.971409449;
cosLookup[2501] <= 0.971386682;
cosLookup[2502] <= 0.971363905;
cosLookup[2503] <= 0.97134112;
cosLookup[2504] <= 0.971318326;
cosLookup[2505] <= 0.971295523;
cosLookup[2506] <= 0.971272711;
cosLookup[2507] <= 0.97124989;
cosLookup[2508] <= 0.971227061;
cosLookup[2509] <= 0.971204222;
cosLookup[2510] <= 0.971181374;
cosLookup[2511] <= 0.971158518;
cosLookup[2512] <= 0.971135652;
cosLookup[2513] <= 0.971112778;
cosLookup[2514] <= 0.971089894;
cosLookup[2515] <= 0.971067002;
cosLookup[2516] <= 0.971044101;
cosLookup[2517] <= 0.971021191;
cosLookup[2518] <= 0.970998272;
cosLookup[2519] <= 0.970975344;
cosLookup[2520] <= 0.970952407;
cosLookup[2521] <= 0.970929461;
cosLookup[2522] <= 0.970906506;
cosLookup[2523] <= 0.970883542;
cosLookup[2524] <= 0.97086057;
cosLookup[2525] <= 0.970837588;
cosLookup[2526] <= 0.970814598;
cosLookup[2527] <= 0.970791598;
cosLookup[2528] <= 0.97076859;
cosLookup[2529] <= 0.970745573;
cosLookup[2530] <= 0.970722547;
cosLookup[2531] <= 0.970699512;
cosLookup[2532] <= 0.970676468;
cosLookup[2533] <= 0.970653415;
cosLookup[2534] <= 0.970630353;
cosLookup[2535] <= 0.970607282;
cosLookup[2536] <= 0.970584202;
cosLookup[2537] <= 0.970561114;
cosLookup[2538] <= 0.970538016;
cosLookup[2539] <= 0.97051491;
cosLookup[2540] <= 0.970491794;
cosLookup[2541] <= 0.97046867;
cosLookup[2542] <= 0.970445537;
cosLookup[2543] <= 0.970422394;
cosLookup[2544] <= 0.970399243;
cosLookup[2545] <= 0.970376083;
cosLookup[2546] <= 0.970352914;
cosLookup[2547] <= 0.970329737;
cosLookup[2548] <= 0.97030655;
cosLookup[2549] <= 0.970283354;
cosLookup[2550] <= 0.97026015;
cosLookup[2551] <= 0.970236936;
cosLookup[2552] <= 0.970213714;
cosLookup[2553] <= 0.970190482;
cosLookup[2554] <= 0.970167242;
cosLookup[2555] <= 0.970143993;
cosLookup[2556] <= 0.970120735;
cosLookup[2557] <= 0.970097468;
cosLookup[2558] <= 0.970074192;
cosLookup[2559] <= 0.970050907;
cosLookup[2560] <= 0.970027613;
cosLookup[2561] <= 0.97000431;
cosLookup[2562] <= 0.969980999;
cosLookup[2563] <= 0.969957678;
cosLookup[2564] <= 0.969934349;
cosLookup[2565] <= 0.96991101;
cosLookup[2566] <= 0.969887663;
cosLookup[2567] <= 0.969864307;
cosLookup[2568] <= 0.969840942;
cosLookup[2569] <= 0.969817568;
cosLookup[2570] <= 0.969794185;
cosLookup[2571] <= 0.969770793;
cosLookup[2572] <= 0.969747392;
cosLookup[2573] <= 0.969723982;
cosLookup[2574] <= 0.969700564;
cosLookup[2575] <= 0.969677136;
cosLookup[2576] <= 0.9696537;
cosLookup[2577] <= 0.969630254;
cosLookup[2578] <= 0.9696068;
cosLookup[2579] <= 0.969583337;
cosLookup[2580] <= 0.969559865;
cosLookup[2581] <= 0.969536384;
cosLookup[2582] <= 0.969512894;
cosLookup[2583] <= 0.969489395;
cosLookup[2584] <= 0.969465887;
cosLookup[2585] <= 0.969442371;
cosLookup[2586] <= 0.969418845;
cosLookup[2587] <= 0.969395311;
cosLookup[2588] <= 0.969371767;
cosLookup[2589] <= 0.969348215;
cosLookup[2590] <= 0.969324654;
cosLookup[2591] <= 0.969301084;
cosLookup[2592] <= 0.969277504;
cosLookup[2593] <= 0.969253917;
cosLookup[2594] <= 0.96923032;
cosLookup[2595] <= 0.969206714;
cosLookup[2596] <= 0.969183099;
cosLookup[2597] <= 0.969159476;
cosLookup[2598] <= 0.969135843;
cosLookup[2599] <= 0.969112202;
cosLookup[2600] <= 0.969088551;
cosLookup[2601] <= 0.969064892;
cosLookup[2602] <= 0.969041224;
cosLookup[2603] <= 0.969017547;
cosLookup[2604] <= 0.968993861;
cosLookup[2605] <= 0.968970166;
cosLookup[2606] <= 0.968946462;
cosLookup[2607] <= 0.96892275;
cosLookup[2608] <= 0.968899028;
cosLookup[2609] <= 0.968875298;
cosLookup[2610] <= 0.968851558;
cosLookup[2611] <= 0.96882781;
cosLookup[2612] <= 0.968804053;
cosLookup[2613] <= 0.968780287;
cosLookup[2614] <= 0.968756512;
cosLookup[2615] <= 0.968732728;
cosLookup[2616] <= 0.968708935;
cosLookup[2617] <= 0.968685133;
cosLookup[2618] <= 0.968661323;
cosLookup[2619] <= 0.968637503;
cosLookup[2620] <= 0.968613675;
cosLookup[2621] <= 0.968589837;
cosLookup[2622] <= 0.968565991;
cosLookup[2623] <= 0.968542136;
cosLookup[2624] <= 0.968518272;
cosLookup[2625] <= 0.968494399;
cosLookup[2626] <= 0.968470517;
cosLookup[2627] <= 0.968446626;
cosLookup[2628] <= 0.968422726;
cosLookup[2629] <= 0.968398818;
cosLookup[2630] <= 0.9683749;
cosLookup[2631] <= 0.968350974;
cosLookup[2632] <= 0.968327039;
cosLookup[2633] <= 0.968303094;
cosLookup[2634] <= 0.968279141;
cosLookup[2635] <= 0.968255179;
cosLookup[2636] <= 0.968231208;
cosLookup[2637] <= 0.968207229;
cosLookup[2638] <= 0.96818324;
cosLookup[2639] <= 0.968159242;
cosLookup[2640] <= 0.968135236;
cosLookup[2641] <= 0.968111221;
cosLookup[2642] <= 0.968087196;
cosLookup[2643] <= 0.968063163;
cosLookup[2644] <= 0.968039121;
cosLookup[2645] <= 0.96801507;
cosLookup[2646] <= 0.96799101;
cosLookup[2647] <= 0.967966941;
cosLookup[2648] <= 0.967942864;
cosLookup[2649] <= 0.967918777;
cosLookup[2650] <= 0.967894681;
cosLookup[2651] <= 0.967870577;
cosLookup[2652] <= 0.967846464;
cosLookup[2653] <= 0.967822342;
cosLookup[2654] <= 0.967798211;
cosLookup[2655] <= 0.967774071;
cosLookup[2656] <= 0.967749922;
cosLookup[2657] <= 0.967725764;
cosLookup[2658] <= 0.967701597;
cosLookup[2659] <= 0.967677422;
cosLookup[2660] <= 0.967653237;
cosLookup[2661] <= 0.967629044;
cosLookup[2662] <= 0.967604842;
cosLookup[2663] <= 0.967580631;
cosLookup[2664] <= 0.967556411;
cosLookup[2665] <= 0.967532182;
cosLookup[2666] <= 0.967507944;
cosLookup[2667] <= 0.967483697;
cosLookup[2668] <= 0.967459441;
cosLookup[2669] <= 0.967435177;
cosLookup[2670] <= 0.967410904;
cosLookup[2671] <= 0.967386621;
cosLookup[2672] <= 0.96736233;
cosLookup[2673] <= 0.96733803;
cosLookup[2674] <= 0.967313721;
cosLookup[2675] <= 0.967289403;
cosLookup[2676] <= 0.967265076;
cosLookup[2677] <= 0.967240741;
cosLookup[2678] <= 0.967216396;
cosLookup[2679] <= 0.967192043;
cosLookup[2680] <= 0.96716768;
cosLookup[2681] <= 0.967143309;
cosLookup[2682] <= 0.967118929;
cosLookup[2683] <= 0.96709454;
cosLookup[2684] <= 0.967070142;
cosLookup[2685] <= 0.967045735;
cosLookup[2686] <= 0.96702132;
cosLookup[2687] <= 0.966996895;
cosLookup[2688] <= 0.966972462;
cosLookup[2689] <= 0.966948019;
cosLookup[2690] <= 0.966923568;
cosLookup[2691] <= 0.966899108;
cosLookup[2692] <= 0.966874639;
cosLookup[2693] <= 0.966850161;
cosLookup[2694] <= 0.966825674;
cosLookup[2695] <= 0.966801179;
cosLookup[2696] <= 0.966776674;
cosLookup[2697] <= 0.966752161;
cosLookup[2698] <= 0.966727639;
cosLookup[2699] <= 0.966703107;
cosLookup[2700] <= 0.966678567;
cosLookup[2701] <= 0.966654018;
cosLookup[2702] <= 0.96662946;
cosLookup[2703] <= 0.966604894;
cosLookup[2704] <= 0.966580318;
cosLookup[2705] <= 0.966555733;
cosLookup[2706] <= 0.96653114;
cosLookup[2707] <= 0.966506538;
cosLookup[2708] <= 0.966481926;
cosLookup[2709] <= 0.966457306;
cosLookup[2710] <= 0.966432677;
cosLookup[2711] <= 0.96640804;
cosLookup[2712] <= 0.966383393;
cosLookup[2713] <= 0.966358737;
cosLookup[2714] <= 0.966334073;
cosLookup[2715] <= 0.966309399;
cosLookup[2716] <= 0.966284717;
cosLookup[2717] <= 0.966260026;
cosLookup[2718] <= 0.966235326;
cosLookup[2719] <= 0.966210617;
cosLookup[2720] <= 0.966185899;
cosLookup[2721] <= 0.966161173;
cosLookup[2722] <= 0.966136437;
cosLookup[2723] <= 0.966111693;
cosLookup[2724] <= 0.966086939;
cosLookup[2725] <= 0.966062177;
cosLookup[2726] <= 0.966037406;
cosLookup[2727] <= 0.966012626;
cosLookup[2728] <= 0.965987837;
cosLookup[2729] <= 0.96596304;
cosLookup[2730] <= 0.965938233;
cosLookup[2731] <= 0.965913417;
cosLookup[2732] <= 0.965888593;
cosLookup[2733] <= 0.96586376;
cosLookup[2734] <= 0.965838918;
cosLookup[2735] <= 0.965814067;
cosLookup[2736] <= 0.965789207;
cosLookup[2737] <= 0.965764338;
cosLookup[2738] <= 0.96573946;
cosLookup[2739] <= 0.965714574;
cosLookup[2740] <= 0.965689679;
cosLookup[2741] <= 0.965664774;
cosLookup[2742] <= 0.965639861;
cosLookup[2743] <= 0.965614939;
cosLookup[2744] <= 0.965590008;
cosLookup[2745] <= 0.965565068;
cosLookup[2746] <= 0.96554012;
cosLookup[2747] <= 0.965515162;
cosLookup[2748] <= 0.965490196;
cosLookup[2749] <= 0.965465221;
cosLookup[2750] <= 0.965440236;
cosLookup[2751] <= 0.965415243;
cosLookup[2752] <= 0.965390242;
cosLookup[2753] <= 0.965365231;
cosLookup[2754] <= 0.965340211;
cosLookup[2755] <= 0.965315183;
cosLookup[2756] <= 0.965290145;
cosLookup[2757] <= 0.965265099;
cosLookup[2758] <= 0.965240044;
cosLookup[2759] <= 0.96521498;
cosLookup[2760] <= 0.965189907;
cosLookup[2761] <= 0.965164825;
cosLookup[2762] <= 0.965139734;
cosLookup[2763] <= 0.965114635;
cosLookup[2764] <= 0.965089527;
cosLookup[2765] <= 0.965064409;
cosLookup[2766] <= 0.965039283;
cosLookup[2767] <= 0.965014148;
cosLookup[2768] <= 0.964989004;
cosLookup[2769] <= 0.964963852;
cosLookup[2770] <= 0.96493869;
cosLookup[2771] <= 0.964913519;
cosLookup[2772] <= 0.96488834;
cosLookup[2773] <= 0.964863152;
cosLookup[2774] <= 0.964837955;
cosLookup[2775] <= 0.964812749;
cosLookup[2776] <= 0.964787534;
cosLookup[2777] <= 0.96476231;
cosLookup[2778] <= 0.964737078;
cosLookup[2779] <= 0.964711836;
cosLookup[2780] <= 0.964686586;
cosLookup[2781] <= 0.964661327;
cosLookup[2782] <= 0.964636059;
cosLookup[2783] <= 0.964610782;
cosLookup[2784] <= 0.964585496;
cosLookup[2785] <= 0.964560201;
cosLookup[2786] <= 0.964534898;
cosLookup[2787] <= 0.964509586;
cosLookup[2788] <= 0.964484264;
cosLookup[2789] <= 0.964458934;
cosLookup[2790] <= 0.964433595;
cosLookup[2791] <= 0.964408247;
cosLookup[2792] <= 0.964382891;
cosLookup[2793] <= 0.964357525;
cosLookup[2794] <= 0.964332151;
cosLookup[2795] <= 0.964306767;
cosLookup[2796] <= 0.964281375;
cosLookup[2797] <= 0.964255974;
cosLookup[2798] <= 0.964230564;
cosLookup[2799] <= 0.964205145;
cosLookup[2800] <= 0.964179718;
cosLookup[2801] <= 0.964154281;
cosLookup[2802] <= 0.964128836;
cosLookup[2803] <= 0.964103382;
cosLookup[2804] <= 0.964077919;
cosLookup[2805] <= 0.964052447;
cosLookup[2806] <= 0.964026966;
cosLookup[2807] <= 0.964001476;
cosLookup[2808] <= 0.963975978;
cosLookup[2809] <= 0.96395047;
cosLookup[2810] <= 0.963924954;
cosLookup[2811] <= 0.963899429;
cosLookup[2812] <= 0.963873895;
cosLookup[2813] <= 0.963848352;
cosLookup[2814] <= 0.9638228;
cosLookup[2815] <= 0.96379724;
cosLookup[2816] <= 0.96377167;
cosLookup[2817] <= 0.963746092;
cosLookup[2818] <= 0.963720505;
cosLookup[2819] <= 0.963694909;
cosLookup[2820] <= 0.963669304;
cosLookup[2821] <= 0.96364369;
cosLookup[2822] <= 0.963618068;
cosLookup[2823] <= 0.963592436;
cosLookup[2824] <= 0.963566796;
cosLookup[2825] <= 0.963541147;
cosLookup[2826] <= 0.963515489;
cosLookup[2827] <= 0.963489822;
cosLookup[2828] <= 0.963464146;
cosLookup[2829] <= 0.963438462;
cosLookup[2830] <= 0.963412768;
cosLookup[2831] <= 0.963387066;
cosLookup[2832] <= 0.963361355;
cosLookup[2833] <= 0.963335635;
cosLookup[2834] <= 0.963309906;
cosLookup[2835] <= 0.963284168;
cosLookup[2836] <= 0.963258422;
cosLookup[2837] <= 0.963232666;
cosLookup[2838] <= 0.963206902;
cosLookup[2839] <= 0.963181129;
cosLookup[2840] <= 0.963155347;
cosLookup[2841] <= 0.963129556;
cosLookup[2842] <= 0.963103756;
cosLookup[2843] <= 0.963077948;
cosLookup[2844] <= 0.96305213;
cosLookup[2845] <= 0.963026304;
cosLookup[2846] <= 0.963000469;
cosLookup[2847] <= 0.962974625;
cosLookup[2848] <= 0.962948772;
cosLookup[2849] <= 0.962922911;
cosLookup[2850] <= 0.96289704;
cosLookup[2851] <= 0.962871161;
cosLookup[2852] <= 0.962845273;
cosLookup[2853] <= 0.962819375;
cosLookup[2854] <= 0.962793469;
cosLookup[2855] <= 0.962767555;
cosLookup[2856] <= 0.962741631;
cosLookup[2857] <= 0.962715699;
cosLookup[2858] <= 0.962689757;
cosLookup[2859] <= 0.962663807;
cosLookup[2860] <= 0.962637848;
cosLookup[2861] <= 0.96261188;
cosLookup[2862] <= 0.962585903;
cosLookup[2863] <= 0.962559918;
cosLookup[2864] <= 0.962533923;
cosLookup[2865] <= 0.96250792;
cosLookup[2866] <= 0.962481908;
cosLookup[2867] <= 0.962455887;
cosLookup[2868] <= 0.962429857;
cosLookup[2869] <= 0.962403819;
cosLookup[2870] <= 0.962377771;
cosLookup[2871] <= 0.962351715;
cosLookup[2872] <= 0.96232565;
cosLookup[2873] <= 0.962299575;
cosLookup[2874] <= 0.962273493;
cosLookup[2875] <= 0.962247401;
cosLookup[2876] <= 0.9622213;
cosLookup[2877] <= 0.962195191;
cosLookup[2878] <= 0.962169073;
cosLookup[2879] <= 0.962142945;
cosLookup[2880] <= 0.962116809;
cosLookup[2881] <= 0.962090665;
cosLookup[2882] <= 0.962064511;
cosLookup[2883] <= 0.962038348;
cosLookup[2884] <= 0.962012177;
cosLookup[2885] <= 0.961985997;
cosLookup[2886] <= 0.961959808;
cosLookup[2887] <= 0.96193361;
cosLookup[2888] <= 0.961907403;
cosLookup[2889] <= 0.961881188;
cosLookup[2890] <= 0.961854963;
cosLookup[2891] <= 0.96182873;
cosLookup[2892] <= 0.961802488;
cosLookup[2893] <= 0.961776237;
cosLookup[2894] <= 0.961749977;
cosLookup[2895] <= 0.961723709;
cosLookup[2896] <= 0.961697431;
cosLookup[2897] <= 0.961671145;
cosLookup[2898] <= 0.96164485;
cosLookup[2899] <= 0.961618546;
cosLookup[2900] <= 0.961592233;
cosLookup[2901] <= 0.961565911;
cosLookup[2902] <= 0.961539581;
cosLookup[2903] <= 0.961513241;
cosLookup[2904] <= 0.961486893;
cosLookup[2905] <= 0.961460536;
cosLookup[2906] <= 0.96143417;
cosLookup[2907] <= 0.961407796;
cosLookup[2908] <= 0.961381412;
cosLookup[2909] <= 0.96135502;
cosLookup[2910] <= 0.961328619;
cosLookup[2911] <= 0.961302209;
cosLookup[2912] <= 0.96127579;
cosLookup[2913] <= 0.961249362;
cosLookup[2914] <= 0.961222925;
cosLookup[2915] <= 0.96119648;
cosLookup[2916] <= 0.961170026;
cosLookup[2917] <= 0.961143563;
cosLookup[2918] <= 0.961117091;
cosLookup[2919] <= 0.96109061;
cosLookup[2920] <= 0.96106412;
cosLookup[2921] <= 0.961037622;
cosLookup[2922] <= 0.961011115;
cosLookup[2923] <= 0.960984599;
cosLookup[2924] <= 0.960958074;
cosLookup[2925] <= 0.96093154;
cosLookup[2926] <= 0.960904998;
cosLookup[2927] <= 0.960878446;
cosLookup[2928] <= 0.960851886;
cosLookup[2929] <= 0.960825317;
cosLookup[2930] <= 0.960798739;
cosLookup[2931] <= 0.960772152;
cosLookup[2932] <= 0.960745557;
cosLookup[2933] <= 0.960718952;
cosLookup[2934] <= 0.960692339;
cosLookup[2935] <= 0.960665717;
cosLookup[2936] <= 0.960639086;
cosLookup[2937] <= 0.960612446;
cosLookup[2938] <= 0.960585798;
cosLookup[2939] <= 0.96055914;
cosLookup[2940] <= 0.960532474;
cosLookup[2941] <= 0.960505799;
cosLookup[2942] <= 0.960479115;
cosLookup[2943] <= 0.960452422;
cosLookup[2944] <= 0.960425721;
cosLookup[2945] <= 0.96039901;
cosLookup[2946] <= 0.960372291;
cosLookup[2947] <= 0.960345563;
cosLookup[2948] <= 0.960318826;
cosLookup[2949] <= 0.960292081;
cosLookup[2950] <= 0.960265326;
cosLookup[2951] <= 0.960238563;
cosLookup[2952] <= 0.960211791;
cosLookup[2953] <= 0.96018501;
cosLookup[2954] <= 0.96015822;
cosLookup[2955] <= 0.960131421;
cosLookup[2956] <= 0.960104614;
cosLookup[2957] <= 0.960077797;
cosLookup[2958] <= 0.960050972;
cosLookup[2959] <= 0.960024138;
cosLookup[2960] <= 0.959997296;
cosLookup[2961] <= 0.959970444;
cosLookup[2962] <= 0.959943584;
cosLookup[2963] <= 0.959916714;
cosLookup[2964] <= 0.959889836;
cosLookup[2965] <= 0.959862949;
cosLookup[2966] <= 0.959836054;
cosLookup[2967] <= 0.959809149;
cosLookup[2968] <= 0.959782236;
cosLookup[2969] <= 0.959755313;
cosLookup[2970] <= 0.959728382;
cosLookup[2971] <= 0.959701443;
cosLookup[2972] <= 0.959674494;
cosLookup[2973] <= 0.959647536;
cosLookup[2974] <= 0.95962057;
cosLookup[2975] <= 0.959593595;
cosLookup[2976] <= 0.959566611;
cosLookup[2977] <= 0.959539618;
cosLookup[2978] <= 0.959512617;
cosLookup[2979] <= 0.959485606;
cosLookup[2980] <= 0.959458587;
cosLookup[2981] <= 0.959431559;
cosLookup[2982] <= 0.959404522;
cosLookup[2983] <= 0.959377476;
cosLookup[2984] <= 0.959350422;
cosLookup[2985] <= 0.959323359;
cosLookup[2986] <= 0.959296286;
cosLookup[2987] <= 0.959269205;
cosLookup[2988] <= 0.959242116;
cosLookup[2989] <= 0.959215017;
cosLookup[2990] <= 0.95918791;
cosLookup[2991] <= 0.959160793;
cosLookup[2992] <= 0.959133668;
cosLookup[2993] <= 0.959106534;
cosLookup[2994] <= 0.959079392;
cosLookup[2995] <= 0.95905224;
cosLookup[2996] <= 0.95902508;
cosLookup[2997] <= 0.958997911;
cosLookup[2998] <= 0.958970733;
cosLookup[2999] <= 0.958943546;
cosLookup[3000] <= 0.95891635;
cosLookup[3001] <= 0.958889146;
cosLookup[3002] <= 0.958861933;
cosLookup[3003] <= 0.958834711;
cosLookup[3004] <= 0.95880748;
cosLookup[3005] <= 0.95878024;
cosLookup[3006] <= 0.958752992;
cosLookup[3007] <= 0.958725734;
cosLookup[3008] <= 0.958698468;
cosLookup[3009] <= 0.958671193;
cosLookup[3010] <= 0.95864391;
cosLookup[3011] <= 0.958616617;
cosLookup[3012] <= 0.958589316;
cosLookup[3013] <= 0.958562006;
cosLookup[3014] <= 0.958534687;
cosLookup[3015] <= 0.958507359;
cosLookup[3016] <= 0.958480022;
cosLookup[3017] <= 0.958452677;
cosLookup[3018] <= 0.958425323;
cosLookup[3019] <= 0.95839796;
cosLookup[3020] <= 0.958370588;
cosLookup[3021] <= 0.958343207;
cosLookup[3022] <= 0.958315818;
cosLookup[3023] <= 0.958288419;
cosLookup[3024] <= 0.958261012;
cosLookup[3025] <= 0.958233596;
cosLookup[3026] <= 0.958206172;
cosLookup[3027] <= 0.958178738;
cosLookup[3028] <= 0.958151296;
cosLookup[3029] <= 0.958123845;
cosLookup[3030] <= 0.958096385;
cosLookup[3031] <= 0.958068916;
cosLookup[3032] <= 0.958041438;
cosLookup[3033] <= 0.958013952;
cosLookup[3034] <= 0.957986457;
cosLookup[3035] <= 0.957958953;
cosLookup[3036] <= 0.95793144;
cosLookup[3037] <= 0.957903919;
cosLookup[3038] <= 0.957876388;
cosLookup[3039] <= 0.957848849;
cosLookup[3040] <= 0.957821301;
cosLookup[3041] <= 0.957793744;
cosLookup[3042] <= 0.957766178;
cosLookup[3043] <= 0.957738604;
cosLookup[3044] <= 0.957711021;
cosLookup[3045] <= 0.957683429;
cosLookup[3046] <= 0.957655828;
cosLookup[3047] <= 0.957628218;
cosLookup[3048] <= 0.9576006;
cosLookup[3049] <= 0.957572973;
cosLookup[3050] <= 0.957545337;
cosLookup[3051] <= 0.957517692;
cosLookup[3052] <= 0.957490038;
cosLookup[3053] <= 0.957462376;
cosLookup[3054] <= 0.957434704;
cosLookup[3055] <= 0.957407024;
cosLookup[3056] <= 0.957379336;
cosLookup[3057] <= 0.957351638;
cosLookup[3058] <= 0.957323931;
cosLookup[3059] <= 0.957296216;
cosLookup[3060] <= 0.957268492;
cosLookup[3061] <= 0.957240759;
cosLookup[3062] <= 0.957213018;
cosLookup[3063] <= 0.957185267;
cosLookup[3064] <= 0.957157508;
cosLookup[3065] <= 0.95712974;
cosLookup[3066] <= 0.957101963;
cosLookup[3067] <= 0.957074177;
cosLookup[3068] <= 0.957046383;
cosLookup[3069] <= 0.95701858;
cosLookup[3070] <= 0.956990767;
cosLookup[3071] <= 0.956962947;
cosLookup[3072] <= 0.956935117;
cosLookup[3073] <= 0.956907279;
cosLookup[3074] <= 0.956879431;
cosLookup[3075] <= 0.956851575;
cosLookup[3076] <= 0.95682371;
cosLookup[3077] <= 0.956795837;
cosLookup[3078] <= 0.956767954;
cosLookup[3079] <= 0.956740063;
cosLookup[3080] <= 0.956712163;
cosLookup[3081] <= 0.956684254;
cosLookup[3082] <= 0.956656337;
cosLookup[3083] <= 0.95662841;
cosLookup[3084] <= 0.956600475;
cosLookup[3085] <= 0.956572531;
cosLookup[3086] <= 0.956544578;
cosLookup[3087] <= 0.956516617;
cosLookup[3088] <= 0.956488646;
cosLookup[3089] <= 0.956460667;
cosLookup[3090] <= 0.956432679;
cosLookup[3091] <= 0.956404683;
cosLookup[3092] <= 0.956376677;
cosLookup[3093] <= 0.956348663;
cosLookup[3094] <= 0.95632064;
cosLookup[3095] <= 0.956292608;
cosLookup[3096] <= 0.956264567;
cosLookup[3097] <= 0.956236518;
cosLookup[3098] <= 0.956208459;
cosLookup[3099] <= 0.956180392;
cosLookup[3100] <= 0.956152316;
cosLookup[3101] <= 0.956124232;
cosLookup[3102] <= 0.956096138;
cosLookup[3103] <= 0.956068036;
cosLookup[3104] <= 0.956039925;
cosLookup[3105] <= 0.956011805;
cosLookup[3106] <= 0.955983677;
cosLookup[3107] <= 0.955955539;
cosLookup[3108] <= 0.955927393;
cosLookup[3109] <= 0.955899238;
cosLookup[3110] <= 0.955871074;
cosLookup[3111] <= 0.955842902;
cosLookup[3112] <= 0.95581472;
cosLookup[3113] <= 0.95578653;
cosLookup[3114] <= 0.955758331;
cosLookup[3115] <= 0.955730124;
cosLookup[3116] <= 0.955701907;
cosLookup[3117] <= 0.955673682;
cosLookup[3118] <= 0.955645448;
cosLookup[3119] <= 0.955617205;
cosLookup[3120] <= 0.955588954;
cosLookup[3121] <= 0.955560693;
cosLookup[3122] <= 0.955532424;
cosLookup[3123] <= 0.955504146;
cosLookup[3124] <= 0.955475859;
cosLookup[3125] <= 0.955447564;
cosLookup[3126] <= 0.955419259;
cosLookup[3127] <= 0.955390946;
cosLookup[3128] <= 0.955362624;
cosLookup[3129] <= 0.955334294;
cosLookup[3130] <= 0.955305954;
cosLookup[3131] <= 0.955277606;
cosLookup[3132] <= 0.955249249;
cosLookup[3133] <= 0.955220883;
cosLookup[3134] <= 0.955192509;
cosLookup[3135] <= 0.955164125;
cosLookup[3136] <= 0.955135733;
cosLookup[3137] <= 0.955107332;
cosLookup[3138] <= 0.955078923;
cosLookup[3139] <= 0.955050504;
cosLookup[3140] <= 0.955022077;
cosLookup[3141] <= 0.954993641;
cosLookup[3142] <= 0.954965196;
cosLookup[3143] <= 0.954936742;
cosLookup[3144] <= 0.95490828;
cosLookup[3145] <= 0.954879809;
cosLookup[3146] <= 0.954851329;
cosLookup[3147] <= 0.95482284;
cosLookup[3148] <= 0.954794343;
cosLookup[3149] <= 0.954765837;
cosLookup[3150] <= 0.954737321;
cosLookup[3151] <= 0.954708798;
cosLookup[3152] <= 0.954680265;
cosLookup[3153] <= 0.954651724;
cosLookup[3154] <= 0.954623174;
cosLookup[3155] <= 0.954594615;
cosLookup[3156] <= 0.954566047;
cosLookup[3157] <= 0.95453747;
cosLookup[3158] <= 0.954508885;
cosLookup[3159] <= 0.954480291;
cosLookup[3160] <= 0.954451688;
cosLookup[3161] <= 0.954423077;
cosLookup[3162] <= 0.954394457;
cosLookup[3163] <= 0.954365827;
cosLookup[3164] <= 0.95433719;
cosLookup[3165] <= 0.954308543;
cosLookup[3166] <= 0.954279887;
cosLookup[3167] <= 0.954251223;
cosLookup[3168] <= 0.95422255;
cosLookup[3169] <= 0.954193868;
cosLookup[3170] <= 0.954165178;
cosLookup[3171] <= 0.954136479;
cosLookup[3172] <= 0.954107771;
cosLookup[3173] <= 0.954079054;
cosLookup[3174] <= 0.954050328;
cosLookup[3175] <= 0.954021594;
cosLookup[3176] <= 0.953992851;
cosLookup[3177] <= 0.953964099;
cosLookup[3178] <= 0.953935338;
cosLookup[3179] <= 0.953906569;
cosLookup[3180] <= 0.95387779;
cosLookup[3181] <= 0.953849003;
cosLookup[3182] <= 0.953820208;
cosLookup[3183] <= 0.953791403;
cosLookup[3184] <= 0.95376259;
cosLookup[3185] <= 0.953733768;
cosLookup[3186] <= 0.953704937;
cosLookup[3187] <= 0.953676097;
cosLookup[3188] <= 0.953647249;
cosLookup[3189] <= 0.953618392;
cosLookup[3190] <= 0.953589526;
cosLookup[3191] <= 0.953560651;
cosLookup[3192] <= 0.953531768;
cosLookup[3193] <= 0.953502876;
cosLookup[3194] <= 0.953473975;
cosLookup[3195] <= 0.953445065;
cosLookup[3196] <= 0.953416146;
cosLookup[3197] <= 0.953387219;
cosLookup[3198] <= 0.953358283;
cosLookup[3199] <= 0.953329338;
cosLookup[3200] <= 0.953300385;
cosLookup[3201] <= 0.953271422;
cosLookup[3202] <= 0.953242451;
cosLookup[3203] <= 0.953213471;
cosLookup[3204] <= 0.953184483;
cosLookup[3205] <= 0.953155485;
cosLookup[3206] <= 0.953126479;
cosLookup[3207] <= 0.953097464;
cosLookup[3208] <= 0.953068441;
cosLookup[3209] <= 0.953039408;
cosLookup[3210] <= 0.953010367;
cosLookup[3211] <= 0.952981317;
cosLookup[3212] <= 0.952952259;
cosLookup[3213] <= 0.952923191;
cosLookup[3214] <= 0.952894115;
cosLookup[3215] <= 0.95286503;
cosLookup[3216] <= 0.952835936;
cosLookup[3217] <= 0.952806834;
cosLookup[3218] <= 0.952777722;
cosLookup[3219] <= 0.952748602;
cosLookup[3220] <= 0.952719474;
cosLookup[3221] <= 0.952690336;
cosLookup[3222] <= 0.95266119;
cosLookup[3223] <= 0.952632035;
cosLookup[3224] <= 0.952602871;
cosLookup[3225] <= 0.952573698;
cosLookup[3226] <= 0.952544517;
cosLookup[3227] <= 0.952515327;
cosLookup[3228] <= 0.952486128;
cosLookup[3229] <= 0.95245692;
cosLookup[3230] <= 0.952427704;
cosLookup[3231] <= 0.952398479;
cosLookup[3232] <= 0.952369245;
cosLookup[3233] <= 0.952340003;
cosLookup[3234] <= 0.952310751;
cosLookup[3235] <= 0.952281491;
cosLookup[3236] <= 0.952252222;
cosLookup[3237] <= 0.952222945;
cosLookup[3238] <= 0.952193658;
cosLookup[3239] <= 0.952164363;
cosLookup[3240] <= 0.952135059;
cosLookup[3241] <= 0.952105747;
cosLookup[3242] <= 0.952076425;
cosLookup[3243] <= 0.952047095;
cosLookup[3244] <= 0.952017756;
cosLookup[3245] <= 0.951988408;
cosLookup[3246] <= 0.951959052;
cosLookup[3247] <= 0.951929687;
cosLookup[3248] <= 0.951900313;
cosLookup[3249] <= 0.95187093;
cosLookup[3250] <= 0.951841539;
cosLookup[3251] <= 0.951812139;
cosLookup[3252] <= 0.95178273;
cosLookup[3253] <= 0.951753312;
cosLookup[3254] <= 0.951723886;
cosLookup[3255] <= 0.951694451;
cosLookup[3256] <= 0.951665007;
cosLookup[3257] <= 0.951635554;
cosLookup[3258] <= 0.951606093;
cosLookup[3259] <= 0.951576623;
cosLookup[3260] <= 0.951547144;
cosLookup[3261] <= 0.951517656;
cosLookup[3262] <= 0.95148816;
cosLookup[3263] <= 0.951458654;
cosLookup[3264] <= 0.951429141;
cosLookup[3265] <= 0.951399618;
cosLookup[3266] <= 0.951370087;
cosLookup[3267] <= 0.951340546;
cosLookup[3268] <= 0.951310998;
cosLookup[3269] <= 0.95128144;
cosLookup[3270] <= 0.951251874;
cosLookup[3271] <= 0.951222298;
cosLookup[3272] <= 0.951192715;
cosLookup[3273] <= 0.951163122;
cosLookup[3274] <= 0.951133521;
cosLookup[3275] <= 0.951103911;
cosLookup[3276] <= 0.951074292;
cosLookup[3277] <= 0.951044664;
cosLookup[3278] <= 0.951015028;
cosLookup[3279] <= 0.950985383;
cosLookup[3280] <= 0.950955729;
cosLookup[3281] <= 0.950926067;
cosLookup[3282] <= 0.950896395;
cosLookup[3283] <= 0.950866715;
cosLookup[3284] <= 0.950837026;
cosLookup[3285] <= 0.950807329;
cosLookup[3286] <= 0.950777623;
cosLookup[3287] <= 0.950747908;
cosLookup[3288] <= 0.950718184;
cosLookup[3289] <= 0.950688452;
cosLookup[3290] <= 0.95065871;
cosLookup[3291] <= 0.95062896;
cosLookup[3292] <= 0.950599202;
cosLookup[3293] <= 0.950569434;
cosLookup[3294] <= 0.950539658;
cosLookup[3295] <= 0.950509873;
cosLookup[3296] <= 0.95048008;
cosLookup[3297] <= 0.950450277;
cosLookup[3298] <= 0.950420466;
cosLookup[3299] <= 0.950390646;
cosLookup[3300] <= 0.950360818;
cosLookup[3301] <= 0.95033098;
cosLookup[3302] <= 0.950301134;
cosLookup[3303] <= 0.95027128;
cosLookup[3304] <= 0.950241416;
cosLookup[3305] <= 0.950211544;
cosLookup[3306] <= 0.950181663;
cosLookup[3307] <= 0.950151773;
cosLookup[3308] <= 0.950121875;
cosLookup[3309] <= 0.950091967;
cosLookup[3310] <= 0.950062051;
cosLookup[3311] <= 0.950032127;
cosLookup[3312] <= 0.950002193;
cosLookup[3313] <= 0.949972251;
cosLookup[3314] <= 0.9499423;
cosLookup[3315] <= 0.949912341;
cosLookup[3316] <= 0.949882372;
cosLookup[3317] <= 0.949852395;
cosLookup[3318] <= 0.949822409;
cosLookup[3319] <= 0.949792415;
cosLookup[3320] <= 0.949762412;
cosLookup[3321] <= 0.9497324;
cosLookup[3322] <= 0.949702379;
cosLookup[3323] <= 0.94967235;
cosLookup[3324] <= 0.949642311;
cosLookup[3325] <= 0.949612264;
cosLookup[3326] <= 0.949582209;
cosLookup[3327] <= 0.949552144;
cosLookup[3328] <= 0.949522071;
cosLookup[3329] <= 0.949491989;
cosLookup[3330] <= 0.949461899;
cosLookup[3331] <= 0.9494318;
cosLookup[3332] <= 0.949401692;
cosLookup[3333] <= 0.949371575;
cosLookup[3334] <= 0.949341449;
cosLookup[3335] <= 0.949311315;
cosLookup[3336] <= 0.949281172;
cosLookup[3337] <= 0.949251021;
cosLookup[3338] <= 0.94922086;
cosLookup[3339] <= 0.949190691;
cosLookup[3340] <= 0.949160513;
cosLookup[3341] <= 0.949130327;
cosLookup[3342] <= 0.949100131;
cosLookup[3343] <= 0.949069927;
cosLookup[3344] <= 0.949039715;
cosLookup[3345] <= 0.949009493;
cosLookup[3346] <= 0.948979263;
cosLookup[3347] <= 0.948949024;
cosLookup[3348] <= 0.948918777;
cosLookup[3349] <= 0.94888852;
cosLookup[3350] <= 0.948858255;
cosLookup[3351] <= 0.948827981;
cosLookup[3352] <= 0.948797699;
cosLookup[3353] <= 0.948767408;
cosLookup[3354] <= 0.948737108;
cosLookup[3355] <= 0.948706799;
cosLookup[3356] <= 0.948676481;
cosLookup[3357] <= 0.948646155;
cosLookup[3358] <= 0.94861582;
cosLookup[3359] <= 0.948585477;
cosLookup[3360] <= 0.948555125;
cosLookup[3361] <= 0.948524764;
cosLookup[3362] <= 0.948494394;
cosLookup[3363] <= 0.948464015;
cosLookup[3364] <= 0.948433628;
cosLookup[3365] <= 0.948403232;
cosLookup[3366] <= 0.948372828;
cosLookup[3367] <= 0.948342414;
cosLookup[3368] <= 0.948311992;
cosLookup[3369] <= 0.948281562;
cosLookup[3370] <= 0.948251122;
cosLookup[3371] <= 0.948220674;
cosLookup[3372] <= 0.948190217;
cosLookup[3373] <= 0.948159751;
cosLookup[3374] <= 0.948129277;
cosLookup[3375] <= 0.948098794;
cosLookup[3376] <= 0.948068302;
cosLookup[3377] <= 0.948037802;
cosLookup[3378] <= 0.948007293;
cosLookup[3379] <= 0.947976775;
cosLookup[3380] <= 0.947946248;
cosLookup[3381] <= 0.947915713;
cosLookup[3382] <= 0.947885169;
cosLookup[3383] <= 0.947854616;
cosLookup[3384] <= 0.947824054;
cosLookup[3385] <= 0.947793484;
cosLookup[3386] <= 0.947762905;
cosLookup[3387] <= 0.947732318;
cosLookup[3388] <= 0.947701721;
cosLookup[3389] <= 0.947671116;
cosLookup[3390] <= 0.947640502;
cosLookup[3391] <= 0.94760988;
cosLookup[3392] <= 0.947579249;
cosLookup[3393] <= 0.947548609;
cosLookup[3394] <= 0.94751796;
cosLookup[3395] <= 0.947487303;
cosLookup[3396] <= 0.947456637;
cosLookup[3397] <= 0.947425962;
cosLookup[3398] <= 0.947395279;
cosLookup[3399] <= 0.947364586;
cosLookup[3400] <= 0.947333886;
cosLookup[3401] <= 0.947303176;
cosLookup[3402] <= 0.947272458;
cosLookup[3403] <= 0.947241731;
cosLookup[3404] <= 0.947210995;
cosLookup[3405] <= 0.947180251;
cosLookup[3406] <= 0.947149497;
cosLookup[3407] <= 0.947118736;
cosLookup[3408] <= 0.947087965;
cosLookup[3409] <= 0.947057186;
cosLookup[3410] <= 0.947026398;
cosLookup[3411] <= 0.946995601;
cosLookup[3412] <= 0.946964796;
cosLookup[3413] <= 0.946933982;
cosLookup[3414] <= 0.946903159;
cosLookup[3415] <= 0.946872328;
cosLookup[3416] <= 0.946841487;
cosLookup[3417] <= 0.946810639;
cosLookup[3418] <= 0.946779781;
cosLookup[3419] <= 0.946748915;
cosLookup[3420] <= 0.94671804;
cosLookup[3421] <= 0.946687156;
cosLookup[3422] <= 0.946656264;
cosLookup[3423] <= 0.946625363;
cosLookup[3424] <= 0.946594453;
cosLookup[3425] <= 0.946563534;
cosLookup[3426] <= 0.946532607;
cosLookup[3427] <= 0.946501671;
cosLookup[3428] <= 0.946470726;
cosLookup[3429] <= 0.946439773;
cosLookup[3430] <= 0.946408811;
cosLookup[3431] <= 0.94637784;
cosLookup[3432] <= 0.946346861;
cosLookup[3433] <= 0.946315873;
cosLookup[3434] <= 0.946284876;
cosLookup[3435] <= 0.946253871;
cosLookup[3436] <= 0.946222856;
cosLookup[3437] <= 0.946191833;
cosLookup[3438] <= 0.946160802;
cosLookup[3439] <= 0.946129762;
cosLookup[3440] <= 0.946098713;
cosLookup[3441] <= 0.946067655;
cosLookup[3442] <= 0.946036588;
cosLookup[3443] <= 0.946005513;
cosLookup[3444] <= 0.94597443;
cosLookup[3445] <= 0.945943337;
cosLookup[3446] <= 0.945912236;
cosLookup[3447] <= 0.945881126;
cosLookup[3448] <= 0.945850007;
cosLookup[3449] <= 0.94581888;
cosLookup[3450] <= 0.945787744;
cosLookup[3451] <= 0.9457566;
cosLookup[3452] <= 0.945725446;
cosLookup[3453] <= 0.945694284;
cosLookup[3454] <= 0.945663113;
cosLookup[3455] <= 0.945631934;
cosLookup[3456] <= 0.945600746;
cosLookup[3457] <= 0.945569549;
cosLookup[3458] <= 0.945538344;
cosLookup[3459] <= 0.945507129;
cosLookup[3460] <= 0.945475906;
cosLookup[3461] <= 0.945444675;
cosLookup[3462] <= 0.945413435;
cosLookup[3463] <= 0.945382186;
cosLookup[3464] <= 0.945350928;
cosLookup[3465] <= 0.945319662;
cosLookup[3466] <= 0.945288387;
cosLookup[3467] <= 0.945257103;
cosLookup[3468] <= 0.94522581;
cosLookup[3469] <= 0.945194509;
cosLookup[3470] <= 0.9451632;
cosLookup[3471] <= 0.945131881;
cosLookup[3472] <= 0.945100554;
cosLookup[3473] <= 0.945069218;
cosLookup[3474] <= 0.945037873;
cosLookup[3475] <= 0.94500652;
cosLookup[3476] <= 0.944975158;
cosLookup[3477] <= 0.944943788;
cosLookup[3478] <= 0.944912408;
cosLookup[3479] <= 0.94488102;
cosLookup[3480] <= 0.944849624;
cosLookup[3481] <= 0.944818218;
cosLookup[3482] <= 0.944786804;
cosLookup[3483] <= 0.944755382;
cosLookup[3484] <= 0.94472395;
cosLookup[3485] <= 0.94469251;
cosLookup[3486] <= 0.944661061;
cosLookup[3487] <= 0.944629604;
cosLookup[3488] <= 0.944598138;
cosLookup[3489] <= 0.944566663;
cosLookup[3490] <= 0.944535179;
cosLookup[3491] <= 0.944503687;
cosLookup[3492] <= 0.944472186;
cosLookup[3493] <= 0.944440677;
cosLookup[3494] <= 0.944409158;
cosLookup[3495] <= 0.944377631;
cosLookup[3496] <= 0.944346096;
cosLookup[3497] <= 0.944314552;
cosLookup[3498] <= 0.944282999;
cosLookup[3499] <= 0.944251437;
cosLookup[3500] <= 0.944219867;
cosLookup[3501] <= 0.944188288;
cosLookup[3502] <= 0.9441567;
cosLookup[3503] <= 0.944125104;
cosLookup[3504] <= 0.944093498;
cosLookup[3505] <= 0.944061885;
cosLookup[3506] <= 0.944030262;
cosLookup[3507] <= 0.943998631;
cosLookup[3508] <= 0.943966991;
cosLookup[3509] <= 0.943935343;
cosLookup[3510] <= 0.943903686;
cosLookup[3511] <= 0.94387202;
cosLookup[3512] <= 0.943840346;
cosLookup[3513] <= 0.943808662;
cosLookup[3514] <= 0.943776971;
cosLookup[3515] <= 0.94374527;
cosLookup[3516] <= 0.943713561;
cosLookup[3517] <= 0.943681843;
cosLookup[3518] <= 0.943650117;
cosLookup[3519] <= 0.943618381;
cosLookup[3520] <= 0.943586637;
cosLookup[3521] <= 0.943554885;
cosLookup[3522] <= 0.943523124;
cosLookup[3523] <= 0.943491354;
cosLookup[3524] <= 0.943459575;
cosLookup[3525] <= 0.943427788;
cosLookup[3526] <= 0.943395992;
cosLookup[3527] <= 0.943364187;
cosLookup[3528] <= 0.943332374;
cosLookup[3529] <= 0.943300552;
cosLookup[3530] <= 0.943268722;
cosLookup[3531] <= 0.943236882;
cosLookup[3532] <= 0.943205034;
cosLookup[3533] <= 0.943173178;
cosLookup[3534] <= 0.943141312;
cosLookup[3535] <= 0.943109438;
cosLookup[3536] <= 0.943077556;
cosLookup[3537] <= 0.943045665;
cosLookup[3538] <= 0.943013765;
cosLookup[3539] <= 0.942981856;
cosLookup[3540] <= 0.942949939;
cosLookup[3541] <= 0.942918013;
cosLookup[3542] <= 0.942886078;
cosLookup[3543] <= 0.942854135;
cosLookup[3544] <= 0.942822183;
cosLookup[3545] <= 0.942790222;
cosLookup[3546] <= 0.942758253;
cosLookup[3547] <= 0.942726275;
cosLookup[3548] <= 0.942694288;
cosLookup[3549] <= 0.942662293;
cosLookup[3550] <= 0.942630289;
cosLookup[3551] <= 0.942598276;
cosLookup[3552] <= 0.942566255;
cosLookup[3553] <= 0.942534225;
cosLookup[3554] <= 0.942502186;
cosLookup[3555] <= 0.942470139;
cosLookup[3556] <= 0.942438083;
cosLookup[3557] <= 0.942406018;
cosLookup[3558] <= 0.942373945;
cosLookup[3559] <= 0.942341863;
cosLookup[3560] <= 0.942309772;
cosLookup[3561] <= 0.942277673;
cosLookup[3562] <= 0.942245565;
cosLookup[3563] <= 0.942213448;
cosLookup[3564] <= 0.942181323;
cosLookup[3565] <= 0.942149189;
cosLookup[3566] <= 0.942117047;
cosLookup[3567] <= 0.942084895;
cosLookup[3568] <= 0.942052735;
cosLookup[3569] <= 0.942020567;
cosLookup[3570] <= 0.94198839;
cosLookup[3571] <= 0.941956204;
cosLookup[3572] <= 0.941924009;
cosLookup[3573] <= 0.941891806;
cosLookup[3574] <= 0.941859594;
cosLookup[3575] <= 0.941827374;
cosLookup[3576] <= 0.941795144;
cosLookup[3577] <= 0.941762907;
cosLookup[3578] <= 0.94173066;
cosLookup[3579] <= 0.941698405;
cosLookup[3580] <= 0.941666141;
cosLookup[3581] <= 0.941633869;
cosLookup[3582] <= 0.941601587;
cosLookup[3583] <= 0.941569298;
cosLookup[3584] <= 0.941536999;
cosLookup[3585] <= 0.941504692;
cosLookup[3586] <= 0.941472376;
cosLookup[3587] <= 0.941440052;
cosLookup[3588] <= 0.941407719;
cosLookup[3589] <= 0.941375377;
cosLookup[3590] <= 0.941343027;
cosLookup[3591] <= 0.941310668;
cosLookup[3592] <= 0.9412783;
cosLookup[3593] <= 0.941245924;
cosLookup[3594] <= 0.941213539;
cosLookup[3595] <= 0.941181145;
cosLookup[3596] <= 0.941148743;
cosLookup[3597] <= 0.941116332;
cosLookup[3598] <= 0.941083912;
cosLookup[3599] <= 0.941051484;
cosLookup[3600] <= 0.941019047;
cosLookup[3601] <= 0.940986602;
cosLookup[3602] <= 0.940954147;
cosLookup[3603] <= 0.940921684;
cosLookup[3604] <= 0.940889213;
cosLookup[3605] <= 0.940856733;
cosLookup[3606] <= 0.940824244;
cosLookup[3607] <= 0.940791747;
cosLookup[3608] <= 0.94075924;
cosLookup[3609] <= 0.940726726;
cosLookup[3610] <= 0.940694202;
cosLookup[3611] <= 0.94066167;
cosLookup[3612] <= 0.94062913;
cosLookup[3613] <= 0.94059658;
cosLookup[3614] <= 0.940564022;
cosLookup[3615] <= 0.940531456;
cosLookup[3616] <= 0.94049888;
cosLookup[3617] <= 0.940466296;
cosLookup[3618] <= 0.940433704;
cosLookup[3619] <= 0.940401103;
cosLookup[3620] <= 0.940368493;
cosLookup[3621] <= 0.940335874;
cosLookup[3622] <= 0.940303247;
cosLookup[3623] <= 0.940270611;
cosLookup[3624] <= 0.940237967;
cosLookup[3625] <= 0.940205314;
cosLookup[3626] <= 0.940172652;
cosLookup[3627] <= 0.940139982;
cosLookup[3628] <= 0.940107303;
cosLookup[3629] <= 0.940074615;
cosLookup[3630] <= 0.940041919;
cosLookup[3631] <= 0.940009214;
cosLookup[3632] <= 0.9399765;
cosLookup[3633] <= 0.939943778;
cosLookup[3634] <= 0.939911047;
cosLookup[3635] <= 0.939878308;
cosLookup[3636] <= 0.93984556;
cosLookup[3637] <= 0.939812803;
cosLookup[3638] <= 0.939780037;
cosLookup[3639] <= 0.939747263;
cosLookup[3640] <= 0.939714481;
cosLookup[3641] <= 0.939681689;
cosLookup[3642] <= 0.939648889;
cosLookup[3643] <= 0.939616081;
cosLookup[3644] <= 0.939583264;
cosLookup[3645] <= 0.939550438;
cosLookup[3646] <= 0.939517603;
cosLookup[3647] <= 0.93948476;
cosLookup[3648] <= 0.939451908;
cosLookup[3649] <= 0.939419048;
cosLookup[3650] <= 0.939386179;
cosLookup[3651] <= 0.939353301;
cosLookup[3652] <= 0.939320415;
cosLookup[3653] <= 0.93928752;
cosLookup[3654] <= 0.939254616;
cosLookup[3655] <= 0.939221704;
cosLookup[3656] <= 0.939188783;
cosLookup[3657] <= 0.939155853;
cosLookup[3658] <= 0.939122915;
cosLookup[3659] <= 0.939089969;
cosLookup[3660] <= 0.939057013;
cosLookup[3661] <= 0.939024049;
cosLookup[3662] <= 0.938991076;
cosLookup[3663] <= 0.938958095;
cosLookup[3664] <= 0.938925105;
cosLookup[3665] <= 0.938892107;
cosLookup[3666] <= 0.938859099;
cosLookup[3667] <= 0.938826084;
cosLookup[3668] <= 0.938793059;
cosLookup[3669] <= 0.938760026;
cosLookup[3670] <= 0.938726984;
cosLookup[3671] <= 0.938693934;
cosLookup[3672] <= 0.938660875;
cosLookup[3673] <= 0.938627807;
cosLookup[3674] <= 0.938594731;
cosLookup[3675] <= 0.938561646;
cosLookup[3676] <= 0.938528553;
cosLookup[3677] <= 0.938495451;
cosLookup[3678] <= 0.93846234;
cosLookup[3679] <= 0.93842922;
cosLookup[3680] <= 0.938396092;
cosLookup[3681] <= 0.938362956;
cosLookup[3682] <= 0.938329811;
cosLookup[3683] <= 0.938296657;
cosLookup[3684] <= 0.938263494;
cosLookup[3685] <= 0.938230323;
cosLookup[3686] <= 0.938197143;
cosLookup[3687] <= 0.938163955;
cosLookup[3688] <= 0.938130758;
cosLookup[3689] <= 0.938097552;
cosLookup[3690] <= 0.938064338;
cosLookup[3691] <= 0.938031115;
cosLookup[3692] <= 0.937997884;
cosLookup[3693] <= 0.937964643;
cosLookup[3694] <= 0.937931395;
cosLookup[3695] <= 0.937898137;
cosLookup[3696] <= 0.937864871;
cosLookup[3697] <= 0.937831597;
cosLookup[3698] <= 0.937798313;
cosLookup[3699] <= 0.937765022;
cosLookup[3700] <= 0.937731721;
cosLookup[3701] <= 0.937698412;
cosLookup[3702] <= 0.937665094;
cosLookup[3703] <= 0.937631768;
cosLookup[3704] <= 0.937598433;
cosLookup[3705] <= 0.937565089;
cosLookup[3706] <= 0.937531737;
cosLookup[3707] <= 0.937498376;
cosLookup[3708] <= 0.937465007;
cosLookup[3709] <= 0.937431629;
cosLookup[3710] <= 0.937398242;
cosLookup[3711] <= 0.937364847;
cosLookup[3712] <= 0.937331443;
cosLookup[3713] <= 0.937298031;
cosLookup[3714] <= 0.937264609;
cosLookup[3715] <= 0.93723118;
cosLookup[3716] <= 0.937197741;
cosLookup[3717] <= 0.937164294;
cosLookup[3718] <= 0.937130839;
cosLookup[3719] <= 0.937097374;
cosLookup[3720] <= 0.937063902;
cosLookup[3721] <= 0.93703042;
cosLookup[3722] <= 0.93699693;
cosLookup[3723] <= 0.936963431;
cosLookup[3724] <= 0.936929924;
cosLookup[3725] <= 0.936896408;
cosLookup[3726] <= 0.936862884;
cosLookup[3727] <= 0.936829351;
cosLookup[3728] <= 0.936795809;
cosLookup[3729] <= 0.936762259;
cosLookup[3730] <= 0.9367287;
cosLookup[3731] <= 0.936695132;
cosLookup[3732] <= 0.936661556;
cosLookup[3733] <= 0.936627971;
cosLookup[3734] <= 0.936594378;
cosLookup[3735] <= 0.936560776;
cosLookup[3736] <= 0.936527165;
cosLookup[3737] <= 0.936493546;
cosLookup[3738] <= 0.936459918;
cosLookup[3739] <= 0.936426281;
cosLookup[3740] <= 0.936392636;
cosLookup[3741] <= 0.936358983;
cosLookup[3742] <= 0.93632532;
cosLookup[3743] <= 0.93629165;
cosLookup[3744] <= 0.93625797;
cosLookup[3745] <= 0.936224282;
cosLookup[3746] <= 0.936190585;
cosLookup[3747] <= 0.93615688;
cosLookup[3748] <= 0.936123166;
cosLookup[3749] <= 0.936089444;
cosLookup[3750] <= 0.936055712;
cosLookup[3751] <= 0.936021973;
cosLookup[3752] <= 0.935988224;
cosLookup[3753] <= 0.935954467;
cosLookup[3754] <= 0.935920702;
cosLookup[3755] <= 0.935886928;
cosLookup[3756] <= 0.935853145;
cosLookup[3757] <= 0.935819354;
cosLookup[3758] <= 0.935785554;
cosLookup[3759] <= 0.935751745;
cosLookup[3760] <= 0.935717928;
cosLookup[3761] <= 0.935684102;
cosLookup[3762] <= 0.935650268;
cosLookup[3763] <= 0.935616425;
cosLookup[3764] <= 0.935582573;
cosLookup[3765] <= 0.935548713;
cosLookup[3766] <= 0.935514844;
cosLookup[3767] <= 0.935480967;
cosLookup[3768] <= 0.935447081;
cosLookup[3769] <= 0.935413186;
cosLookup[3770] <= 0.935379283;
cosLookup[3771] <= 0.935345371;
cosLookup[3772] <= 0.935311451;
cosLookup[3773] <= 0.935277522;
cosLookup[3774] <= 0.935243585;
cosLookup[3775] <= 0.935209638;
cosLookup[3776] <= 0.935175684;
cosLookup[3777] <= 0.93514172;
cosLookup[3778] <= 0.935107748;
cosLookup[3779] <= 0.935073768;
cosLookup[3780] <= 0.935039779;
cosLookup[3781] <= 0.935005781;
cosLookup[3782] <= 0.934971775;
cosLookup[3783] <= 0.93493776;
cosLookup[3784] <= 0.934903736;
cosLookup[3785] <= 0.934869704;
cosLookup[3786] <= 0.934835663;
cosLookup[3787] <= 0.934801614;
cosLookup[3788] <= 0.934767556;
cosLookup[3789] <= 0.93473349;
cosLookup[3790] <= 0.934699415;
cosLookup[3791] <= 0.934665331;
cosLookup[3792] <= 0.934631239;
cosLookup[3793] <= 0.934597138;
cosLookup[3794] <= 0.934563028;
cosLookup[3795] <= 0.93452891;
cosLookup[3796] <= 0.934494784;
cosLookup[3797] <= 0.934460648;
cosLookup[3798] <= 0.934426505;
cosLookup[3799] <= 0.934392352;
cosLookup[3800] <= 0.934358191;
cosLookup[3801] <= 0.934324022;
cosLookup[3802] <= 0.934289843;
cosLookup[3803] <= 0.934255657;
cosLookup[3804] <= 0.934221461;
cosLookup[3805] <= 0.934187257;
cosLookup[3806] <= 0.934153045;
cosLookup[3807] <= 0.934118824;
cosLookup[3808] <= 0.934084594;
cosLookup[3809] <= 0.934050356;
cosLookup[3810] <= 0.934016109;
cosLookup[3811] <= 0.933981853;
cosLookup[3812] <= 0.933947589;
cosLookup[3813] <= 0.933913317;
cosLookup[3814] <= 0.933879035;
cosLookup[3815] <= 0.933844746;
cosLookup[3816] <= 0.933810447;
cosLookup[3817] <= 0.93377614;
cosLookup[3818] <= 0.933741825;
cosLookup[3819] <= 0.9337075;
cosLookup[3820] <= 0.933673168;
cosLookup[3821] <= 0.933638826;
cosLookup[3822] <= 0.933604477;
cosLookup[3823] <= 0.933570118;
cosLookup[3824] <= 0.933535751;
cosLookup[3825] <= 0.933501375;
cosLookup[3826] <= 0.933466991;
cosLookup[3827] <= 0.933432598;
cosLookup[3828] <= 0.933398197;
cosLookup[3829] <= 0.933363787;
cosLookup[3830] <= 0.933329368;
cosLookup[3831] <= 0.933294941;
cosLookup[3832] <= 0.933260506;
cosLookup[3833] <= 0.933226061;
cosLookup[3834] <= 0.933191608;
cosLookup[3835] <= 0.933157147;
cosLookup[3836] <= 0.933122677;
cosLookup[3837] <= 0.933088198;
cosLookup[3838] <= 0.933053711;
cosLookup[3839] <= 0.933019215;
cosLookup[3840] <= 0.932984711;
cosLookup[3841] <= 0.932950198;
cosLookup[3842] <= 0.932915677;
cosLookup[3843] <= 0.932881147;
cosLookup[3844] <= 0.932846608;
cosLookup[3845] <= 0.932812061;
cosLookup[3846] <= 0.932777505;
cosLookup[3847] <= 0.932742941;
cosLookup[3848] <= 0.932708368;
cosLookup[3849] <= 0.932673786;
cosLookup[3850] <= 0.932639196;
cosLookup[3851] <= 0.932604597;
cosLookup[3852] <= 0.93256999;
cosLookup[3853] <= 0.932535374;
cosLookup[3854] <= 0.93250075;
cosLookup[3855] <= 0.932466117;
cosLookup[3856] <= 0.932431476;
cosLookup[3857] <= 0.932396825;
cosLookup[3858] <= 0.932362167;
cosLookup[3859] <= 0.9323275;
cosLookup[3860] <= 0.932292824;
cosLookup[3861] <= 0.932258139;
cosLookup[3862] <= 0.932223446;
cosLookup[3863] <= 0.932188745;
cosLookup[3864] <= 0.932154035;
cosLookup[3865] <= 0.932119316;
cosLookup[3866] <= 0.932084589;
cosLookup[3867] <= 0.932049853;
cosLookup[3868] <= 0.932015109;
cosLookup[3869] <= 0.931980356;
cosLookup[3870] <= 0.931945594;
cosLookup[3871] <= 0.931910824;
cosLookup[3872] <= 0.931876046;
cosLookup[3873] <= 0.931841258;
cosLookup[3874] <= 0.931806463;
cosLookup[3875] <= 0.931771658;
cosLookup[3876] <= 0.931736845;
cosLookup[3877] <= 0.931702024;
cosLookup[3878] <= 0.931667194;
cosLookup[3879] <= 0.931632355;
cosLookup[3880] <= 0.931597508;
cosLookup[3881] <= 0.931562652;
cosLookup[3882] <= 0.931527788;
cosLookup[3883] <= 0.931492915;
cosLookup[3884] <= 0.931458034;
cosLookup[3885] <= 0.931423144;
cosLookup[3886] <= 0.931388245;
cosLookup[3887] <= 0.931353338;
cosLookup[3888] <= 0.931318423;
cosLookup[3889] <= 0.931283498;
cosLookup[3890] <= 0.931248566;
cosLookup[3891] <= 0.931213624;
cosLookup[3892] <= 0.931178674;
cosLookup[3893] <= 0.931143716;
cosLookup[3894] <= 0.931108749;
cosLookup[3895] <= 0.931073773;
cosLookup[3896] <= 0.931038789;
cosLookup[3897] <= 0.931003796;
cosLookup[3898] <= 0.930968795;
cosLookup[3899] <= 0.930933785;
cosLookup[3900] <= 0.930898767;
cosLookup[3901] <= 0.93086374;
cosLookup[3902] <= 0.930828705;
cosLookup[3903] <= 0.930793661;
cosLookup[3904] <= 0.930758608;
cosLookup[3905] <= 0.930723547;
cosLookup[3906] <= 0.930688477;
cosLookup[3907] <= 0.930653399;
cosLookup[3908] <= 0.930618312;
cosLookup[3909] <= 0.930583217;
cosLookup[3910] <= 0.930548113;
cosLookup[3911] <= 0.930513;
cosLookup[3912] <= 0.930477879;
cosLookup[3913] <= 0.930442749;
cosLookup[3914] <= 0.930407611;
cosLookup[3915] <= 0.930372465;
cosLookup[3916] <= 0.930337309;
cosLookup[3917] <= 0.930302146;
cosLookup[3918] <= 0.930266973;
cosLookup[3919] <= 0.930231792;
cosLookup[3920] <= 0.930196603;
cosLookup[3921] <= 0.930161405;
cosLookup[3922] <= 0.930126198;
cosLookup[3923] <= 0.930090983;
cosLookup[3924] <= 0.930055759;
cosLookup[3925] <= 0.930020527;
cosLookup[3926] <= 0.929985286;
cosLookup[3927] <= 0.929950037;
cosLookup[3928] <= 0.929914779;
cosLookup[3929] <= 0.929879513;
cosLookup[3930] <= 0.929844238;
cosLookup[3931] <= 0.929808954;
cosLookup[3932] <= 0.929773662;
cosLookup[3933] <= 0.929738362;
cosLookup[3934] <= 0.929703052;
cosLookup[3935] <= 0.929667735;
cosLookup[3936] <= 0.929632408;
cosLookup[3937] <= 0.929597074;
cosLookup[3938] <= 0.92956173;
cosLookup[3939] <= 0.929526378;
cosLookup[3940] <= 0.929491018;
cosLookup[3941] <= 0.929455649;
cosLookup[3942] <= 0.929420272;
cosLookup[3943] <= 0.929384885;
cosLookup[3944] <= 0.929349491;
cosLookup[3945] <= 0.929314088;
cosLookup[3946] <= 0.929278676;
cosLookup[3947] <= 0.929243256;
cosLookup[3948] <= 0.929207827;
cosLookup[3949] <= 0.92917239;
cosLookup[3950] <= 0.929136944;
cosLookup[3951] <= 0.929101489;
cosLookup[3952] <= 0.929066026;
cosLookup[3953] <= 0.929030555;
cosLookup[3954] <= 0.928995075;
cosLookup[3955] <= 0.928959586;
cosLookup[3956] <= 0.928924089;
cosLookup[3957] <= 0.928888584;
cosLookup[3958] <= 0.928853069;
cosLookup[3959] <= 0.928817547;
cosLookup[3960] <= 0.928782015;
cosLookup[3961] <= 0.928746476;
cosLookup[3962] <= 0.928710927;
cosLookup[3963] <= 0.92867537;
cosLookup[3964] <= 0.928639805;
cosLookup[3965] <= 0.928604231;
cosLookup[3966] <= 0.928568649;
cosLookup[3967] <= 0.928533057;
cosLookup[3968] <= 0.928497458;
cosLookup[3969] <= 0.92846185;
cosLookup[3970] <= 0.928426233;
cosLookup[3971] <= 0.928390608;
cosLookup[3972] <= 0.928354974;
cosLookup[3973] <= 0.928319332;
cosLookup[3974] <= 0.928283681;
cosLookup[3975] <= 0.928248022;
cosLookup[3976] <= 0.928212354;
cosLookup[3977] <= 0.928176678;
cosLookup[3978] <= 0.928140993;
cosLookup[3979] <= 0.928105299;
cosLookup[3980] <= 0.928069597;
cosLookup[3981] <= 0.928033887;
cosLookup[3982] <= 0.927998168;
cosLookup[3983] <= 0.92796244;
cosLookup[3984] <= 0.927926704;
cosLookup[3985] <= 0.92789096;
cosLookup[3986] <= 0.927855207;
cosLookup[3987] <= 0.927819445;
cosLookup[3988] <= 0.927783675;
cosLookup[3989] <= 0.927747896;
cosLookup[3990] <= 0.927712109;
cosLookup[3991] <= 0.927676313;
cosLookup[3992] <= 0.927640508;
cosLookup[3993] <= 0.927604696;
cosLookup[3994] <= 0.927568874;
cosLookup[3995] <= 0.927533044;
cosLookup[3996] <= 0.927497206;
cosLookup[3997] <= 0.927461359;
cosLookup[3998] <= 0.927425503;
cosLookup[3999] <= 0.927389639;
cosLookup[4000] <= 0.927353767;
cosLookup[4001] <= 0.927317886;
cosLookup[4002] <= 0.927281996;
cosLookup[4003] <= 0.927246098;
cosLookup[4004] <= 0.927210192;
cosLookup[4005] <= 0.927174276;
cosLookup[4006] <= 0.927138353;
cosLookup[4007] <= 0.92710242;
cosLookup[4008] <= 0.92706648;
cosLookup[4009] <= 0.92703053;
cosLookup[4010] <= 0.926994573;
cosLookup[4011] <= 0.926958606;
cosLookup[4012] <= 0.926922632;
cosLookup[4013] <= 0.926886648;
cosLookup[4014] <= 0.926850656;
cosLookup[4015] <= 0.926814656;
cosLookup[4016] <= 0.926778647;
cosLookup[4017] <= 0.92674263;
cosLookup[4018] <= 0.926706604;
cosLookup[4019] <= 0.926670569;
cosLookup[4020] <= 0.926634526;
cosLookup[4021] <= 0.926598475;
cosLookup[4022] <= 0.926562415;
cosLookup[4023] <= 0.926526346;
cosLookup[4024] <= 0.926490269;
cosLookup[4025] <= 0.926454184;
cosLookup[4026] <= 0.92641809;
cosLookup[4027] <= 0.926381987;
cosLookup[4028] <= 0.926345876;
cosLookup[4029] <= 0.926309756;
cosLookup[4030] <= 0.926273628;
cosLookup[4031] <= 0.926237491;
cosLookup[4032] <= 0.926201346;
cosLookup[4033] <= 0.926165193;
cosLookup[4034] <= 0.92612903;
cosLookup[4035] <= 0.92609286;
cosLookup[4036] <= 0.92605668;
cosLookup[4037] <= 0.926020493;
cosLookup[4038] <= 0.925984296;
cosLookup[4039] <= 0.925948092;
cosLookup[4040] <= 0.925911878;
cosLookup[4041] <= 0.925875657;
cosLookup[4042] <= 0.925839426;
cosLookup[4043] <= 0.925803187;
cosLookup[4044] <= 0.92576694;
cosLookup[4045] <= 0.925730684;
cosLookup[4046] <= 0.92569442;
cosLookup[4047] <= 0.925658147;
cosLookup[4048] <= 0.925621866;
cosLookup[4049] <= 0.925585576;
cosLookup[4050] <= 0.925549277;
cosLookup[4051] <= 0.925512971;
cosLookup[4052] <= 0.925476655;
cosLookup[4053] <= 0.925440331;
cosLookup[4054] <= 0.925403999;
cosLookup[4055] <= 0.925367658;
cosLookup[4056] <= 0.925331308;
cosLookup[4057] <= 0.92529495;
cosLookup[4058] <= 0.925258584;
cosLookup[4059] <= 0.925222209;
cosLookup[4060] <= 0.925185826;
cosLookup[4061] <= 0.925149434;
cosLookup[4062] <= 0.925113033;
cosLookup[4063] <= 0.925076624;
cosLookup[4064] <= 0.925040207;
cosLookup[4065] <= 0.925003781;
cosLookup[4066] <= 0.924967346;
cosLookup[4067] <= 0.924930903;
cosLookup[4068] <= 0.924894452;
cosLookup[4069] <= 0.924857992;
cosLookup[4070] <= 0.924821523;
cosLookup[4071] <= 0.924785046;
cosLookup[4072] <= 0.924748561;
cosLookup[4073] <= 0.924712067;
cosLookup[4074] <= 0.924675564;
cosLookup[4075] <= 0.924639053;
cosLookup[4076] <= 0.924602534;
cosLookup[4077] <= 0.924566006;
cosLookup[4078] <= 0.924529469;
cosLookup[4079] <= 0.924492924;
cosLookup[4080] <= 0.924456371;
cosLookup[4081] <= 0.924419809;
cosLookup[4082] <= 0.924383238;
cosLookup[4083] <= 0.924346659;
cosLookup[4084] <= 0.924310072;
cosLookup[4085] <= 0.924273476;
cosLookup[4086] <= 0.924236871;
cosLookup[4087] <= 0.924200258;
cosLookup[4088] <= 0.924163637;
cosLookup[4089] <= 0.924127007;
cosLookup[4090] <= 0.924090369;
cosLookup[4091] <= 0.924053722;
cosLookup[4092] <= 0.924017066;
cosLookup[4093] <= 0.923980402;
cosLookup[4094] <= 0.92394373;
cosLookup[4095] <= 0.923907049;
cosLookup[4096] <= 0.923870359;
cosLookup[4097] <= 0.923833661;
cosLookup[4098] <= 0.923796955;
cosLookup[4099] <= 0.92376024;
cosLookup[4100] <= 0.923723517;
cosLookup[4101] <= 0.923686785;
cosLookup[4102] <= 0.923650044;
cosLookup[4103] <= 0.923613296;
cosLookup[4104] <= 0.923576538;
cosLookup[4105] <= 0.923539772;
cosLookup[4106] <= 0.923502998;
cosLookup[4107] <= 0.923466215;
cosLookup[4108] <= 0.923429424;
cosLookup[4109] <= 0.923392624;
cosLookup[4110] <= 0.923355816;
cosLookup[4111] <= 0.923318999;
cosLookup[4112] <= 0.923282174;
cosLookup[4113] <= 0.92324534;
cosLookup[4114] <= 0.923208498;
cosLookup[4115] <= 0.923171647;
cosLookup[4116] <= 0.923134788;
cosLookup[4117] <= 0.92309792;
cosLookup[4118] <= 0.923061044;
cosLookup[4119] <= 0.923024159;
cosLookup[4120] <= 0.922987266;
cosLookup[4121] <= 0.922950364;
cosLookup[4122] <= 0.922913454;
cosLookup[4123] <= 0.922876535;
cosLookup[4124] <= 0.922839608;
cosLookup[4125] <= 0.922802673;
cosLookup[4126] <= 0.922765729;
cosLookup[4127] <= 0.922728776;
cosLookup[4128] <= 0.922691815;
cosLookup[4129] <= 0.922654846;
cosLookup[4130] <= 0.922617868;
cosLookup[4131] <= 0.922580881;
cosLookup[4132] <= 0.922543886;
cosLookup[4133] <= 0.922506883;
cosLookup[4134] <= 0.922469871;
cosLookup[4135] <= 0.92243285;
cosLookup[4136] <= 0.922395821;
cosLookup[4137] <= 0.922358784;
cosLookup[4138] <= 0.922321738;
cosLookup[4139] <= 0.922284684;
cosLookup[4140] <= 0.922247621;
cosLookup[4141] <= 0.92221055;
cosLookup[4142] <= 0.92217347;
cosLookup[4143] <= 0.922136382;
cosLookup[4144] <= 0.922099285;
cosLookup[4145] <= 0.92206218;
cosLookup[4146] <= 0.922025066;
cosLookup[4147] <= 0.921987944;
cosLookup[4148] <= 0.921950813;
cosLookup[4149] <= 0.921913674;
cosLookup[4150] <= 0.921876527;
cosLookup[4151] <= 0.921839371;
cosLookup[4152] <= 0.921802206;
cosLookup[4153] <= 0.921765033;
cosLookup[4154] <= 0.921727852;
cosLookup[4155] <= 0.921690662;
cosLookup[4156] <= 0.921653463;
cosLookup[4157] <= 0.921616257;
cosLookup[4158] <= 0.921579041;
cosLookup[4159] <= 0.921541817;
cosLookup[4160] <= 0.921504585;
cosLookup[4161] <= 0.921467344;
cosLookup[4162] <= 0.921430095;
cosLookup[4163] <= 0.921392837;
cosLookup[4164] <= 0.921355571;
cosLookup[4165] <= 0.921318296;
cosLookup[4166] <= 0.921281013;
cosLookup[4167] <= 0.921243722;
cosLookup[4168] <= 0.921206422;
cosLookup[4169] <= 0.921169113;
cosLookup[4170] <= 0.921131796;
cosLookup[4171] <= 0.921094471;
cosLookup[4172] <= 0.921057137;
cosLookup[4173] <= 0.921019794;
cosLookup[4174] <= 0.920982443;
cosLookup[4175] <= 0.920945084;
cosLookup[4176] <= 0.920907716;
cosLookup[4177] <= 0.92087034;
cosLookup[4178] <= 0.920832955;
cosLookup[4179] <= 0.920795562;
cosLookup[4180] <= 0.92075816;
cosLookup[4181] <= 0.92072075;
cosLookup[4182] <= 0.920683332;
cosLookup[4183] <= 0.920645905;
cosLookup[4184] <= 0.920608469;
cosLookup[4185] <= 0.920571025;
cosLookup[4186] <= 0.920533573;
cosLookup[4187] <= 0.920496112;
cosLookup[4188] <= 0.920458642;
cosLookup[4189] <= 0.920421165;
cosLookup[4190] <= 0.920383678;
cosLookup[4191] <= 0.920346184;
cosLookup[4192] <= 0.92030868;
cosLookup[4193] <= 0.920271169;
cosLookup[4194] <= 0.920233649;
cosLookup[4195] <= 0.92019612;
cosLookup[4196] <= 0.920158583;
cosLookup[4197] <= 0.920121037;
cosLookup[4198] <= 0.920083483;
cosLookup[4199] <= 0.920045921;
cosLookup[4200] <= 0.92000835;
cosLookup[4201] <= 0.919970771;
cosLookup[4202] <= 0.919933183;
cosLookup[4203] <= 0.919895587;
cosLookup[4204] <= 0.919857982;
cosLookup[4205] <= 0.919820369;
cosLookup[4206] <= 0.919782747;
cosLookup[4207] <= 0.919745117;
cosLookup[4208] <= 0.919707479;
cosLookup[4209] <= 0.919669832;
cosLookup[4210] <= 0.919632176;
cosLookup[4211] <= 0.919594512;
cosLookup[4212] <= 0.91955684;
cosLookup[4213] <= 0.919519159;
cosLookup[4214] <= 0.91948147;
cosLookup[4215] <= 0.919443772;
cosLookup[4216] <= 0.919406066;
cosLookup[4217] <= 0.919368351;
cosLookup[4218] <= 0.919330628;
cosLookup[4219] <= 0.919292897;
cosLookup[4220] <= 0.919255157;
cosLookup[4221] <= 0.919217408;
cosLookup[4222] <= 0.919179651;
cosLookup[4223] <= 0.919141886;
cosLookup[4224] <= 0.919104112;
cosLookup[4225] <= 0.91906633;
cosLookup[4226] <= 0.919028539;
cosLookup[4227] <= 0.91899074;
cosLookup[4228] <= 0.918952933;
cosLookup[4229] <= 0.918915117;
cosLookup[4230] <= 0.918877292;
cosLookup[4231] <= 0.918839459;
cosLookup[4232] <= 0.918801618;
cosLookup[4233] <= 0.918763768;
cosLookup[4234] <= 0.91872591;
cosLookup[4235] <= 0.918688043;
cosLookup[4236] <= 0.918650168;
cosLookup[4237] <= 0.918612285;
cosLookup[4238] <= 0.918574392;
cosLookup[4239] <= 0.918536492;
cosLookup[4240] <= 0.918498583;
cosLookup[4241] <= 0.918460666;
cosLookup[4242] <= 0.91842274;
cosLookup[4243] <= 0.918384806;
cosLookup[4244] <= 0.918346863;
cosLookup[4245] <= 0.918308912;
cosLookup[4246] <= 0.918270952;
cosLookup[4247] <= 0.918232984;
cosLookup[4248] <= 0.918195008;
cosLookup[4249] <= 0.918157023;
cosLookup[4250] <= 0.91811903;
cosLookup[4251] <= 0.918081028;
cosLookup[4252] <= 0.918043018;
cosLookup[4253] <= 0.918004999;
cosLookup[4254] <= 0.917966972;
cosLookup[4255] <= 0.917928936;
cosLookup[4256] <= 0.917890892;
cosLookup[4257] <= 0.91785284;
cosLookup[4258] <= 0.917814779;
cosLookup[4259] <= 0.91777671;
cosLookup[4260] <= 0.917738632;
cosLookup[4261] <= 0.917700546;
cosLookup[4262] <= 0.917662451;
cosLookup[4263] <= 0.917624348;
cosLookup[4264] <= 0.917586237;
cosLookup[4265] <= 0.917548117;
cosLookup[4266] <= 0.917509988;
cosLookup[4267] <= 0.917471852;
cosLookup[4268] <= 0.917433707;
cosLookup[4269] <= 0.917395553;
cosLookup[4270] <= 0.917357391;
cosLookup[4271] <= 0.91731922;
cosLookup[4272] <= 0.917281041;
cosLookup[4273] <= 0.917242854;
cosLookup[4274] <= 0.917204658;
cosLookup[4275] <= 0.917166454;
cosLookup[4276] <= 0.917128241;
cosLookup[4277] <= 0.91709002;
cosLookup[4278] <= 0.917051791;
cosLookup[4279] <= 0.917013553;
cosLookup[4280] <= 0.916975306;
cosLookup[4281] <= 0.916937051;
cosLookup[4282] <= 0.916898788;
cosLookup[4283] <= 0.916860516;
cosLookup[4284] <= 0.916822236;
cosLookup[4285] <= 0.916783948;
cosLookup[4286] <= 0.916745651;
cosLookup[4287] <= 0.916707345;
cosLookup[4288] <= 0.916669032;
cosLookup[4289] <= 0.916630709;
cosLookup[4290] <= 0.916592379;
cosLookup[4291] <= 0.91655404;
cosLookup[4292] <= 0.916515692;
cosLookup[4293] <= 0.916477336;
cosLookup[4294] <= 0.916438972;
cosLookup[4295] <= 0.916400599;
cosLookup[4296] <= 0.916362218;
cosLookup[4297] <= 0.916323828;
cosLookup[4298] <= 0.91628543;
cosLookup[4299] <= 0.916247024;
cosLookup[4300] <= 0.916208609;
cosLookup[4301] <= 0.916170185;
cosLookup[4302] <= 0.916131754;
cosLookup[4303] <= 0.916093313;
cosLookup[4304] <= 0.916054865;
cosLookup[4305] <= 0.916016408;
cosLookup[4306] <= 0.915977942;
cosLookup[4307] <= 0.915939468;
cosLookup[4308] <= 0.915900986;
cosLookup[4309] <= 0.915862495;
cosLookup[4310] <= 0.915823996;
cosLookup[4311] <= 0.915785489;
cosLookup[4312] <= 0.915746973;
cosLookup[4313] <= 0.915708448;
cosLookup[4314] <= 0.915669916;
cosLookup[4315] <= 0.915631374;
cosLookup[4316] <= 0.915592825;
cosLookup[4317] <= 0.915554267;
cosLookup[4318] <= 0.9155157;
cosLookup[4319] <= 0.915477125;
cosLookup[4320] <= 0.915438542;
cosLookup[4321] <= 0.91539995;
cosLookup[4322] <= 0.91536135;
cosLookup[4323] <= 0.915322742;
cosLookup[4324] <= 0.915284125;
cosLookup[4325] <= 0.915245499;
cosLookup[4326] <= 0.915206865;
cosLookup[4327] <= 0.915168223;
cosLookup[4328] <= 0.915129573;
cosLookup[4329] <= 0.915090914;
cosLookup[4330] <= 0.915052246;
cosLookup[4331] <= 0.91501357;
cosLookup[4332] <= 0.914974886;
cosLookup[4333] <= 0.914936193;
cosLookup[4334] <= 0.914897492;
cosLookup[4335] <= 0.914858783;
cosLookup[4336] <= 0.914820065;
cosLookup[4337] <= 0.914781338;
cosLookup[4338] <= 0.914742604;
cosLookup[4339] <= 0.914703861;
cosLookup[4340] <= 0.914665109;
cosLookup[4341] <= 0.914626349;
cosLookup[4342] <= 0.914587581;
cosLookup[4343] <= 0.914548804;
cosLookup[4344] <= 0.914510019;
cosLookup[4345] <= 0.914471225;
cosLookup[4346] <= 0.914432423;
cosLookup[4347] <= 0.914393613;
cosLookup[4348] <= 0.914354794;
cosLookup[4349] <= 0.914315967;
cosLookup[4350] <= 0.914277131;
cosLookup[4351] <= 0.914238287;
cosLookup[4352] <= 0.914199435;
cosLookup[4353] <= 0.914160574;
cosLookup[4354] <= 0.914121705;
cosLookup[4355] <= 0.914082827;
cosLookup[4356] <= 0.914043941;
cosLookup[4357] <= 0.914005047;
cosLookup[4358] <= 0.913966144;
cosLookup[4359] <= 0.913927232;
cosLookup[4360] <= 0.913888313;
cosLookup[4361] <= 0.913849385;
cosLookup[4362] <= 0.913810448;
cosLookup[4363] <= 0.913771503;
cosLookup[4364] <= 0.91373255;
cosLookup[4365] <= 0.913693589;
cosLookup[4366] <= 0.913654618;
cosLookup[4367] <= 0.91361564;
cosLookup[4368] <= 0.913576653;
cosLookup[4369] <= 0.913537658;
cosLookup[4370] <= 0.913498654;
cosLookup[4371] <= 0.913459642;
cosLookup[4372] <= 0.913420622;
cosLookup[4373] <= 0.913381593;
cosLookup[4374] <= 0.913342556;
cosLookup[4375] <= 0.91330351;
cosLookup[4376] <= 0.913264456;
cosLookup[4377] <= 0.913225394;
cosLookup[4378] <= 0.913186323;
cosLookup[4379] <= 0.913147244;
cosLookup[4380] <= 0.913108156;
cosLookup[4381] <= 0.91306906;
cosLookup[4382] <= 0.913029956;
cosLookup[4383] <= 0.912990843;
cosLookup[4384] <= 0.912951722;
cosLookup[4385] <= 0.912912592;
cosLookup[4386] <= 0.912873454;
cosLookup[4387] <= 0.912834308;
cosLookup[4388] <= 0.912795153;
cosLookup[4389] <= 0.91275599;
cosLookup[4390] <= 0.912716818;
cosLookup[4391] <= 0.912677638;
cosLookup[4392] <= 0.91263845;
cosLookup[4393] <= 0.912599253;
cosLookup[4394] <= 0.912560048;
cosLookup[4395] <= 0.912520835;
cosLookup[4396] <= 0.912481613;
cosLookup[4397] <= 0.912442383;
cosLookup[4398] <= 0.912403144;
cosLookup[4399] <= 0.912363897;
cosLookup[4400] <= 0.912324642;
cosLookup[4401] <= 0.912285378;
cosLookup[4402] <= 0.912246106;
cosLookup[4403] <= 0.912206825;
cosLookup[4404] <= 0.912167536;
cosLookup[4405] <= 0.912128239;
cosLookup[4406] <= 0.912088933;
cosLookup[4407] <= 0.912049619;
cosLookup[4408] <= 0.912010296;
cosLookup[4409] <= 0.911970965;
cosLookup[4410] <= 0.911931626;
cosLookup[4411] <= 0.911892278;
cosLookup[4412] <= 0.911852922;
cosLookup[4413] <= 0.911813558;
cosLookup[4414] <= 0.911774185;
cosLookup[4415] <= 0.911734804;
cosLookup[4416] <= 0.911695414;
cosLookup[4417] <= 0.911656017;
cosLookup[4418] <= 0.91161661;
cosLookup[4419] <= 0.911577195;
cosLookup[4420] <= 0.911537772;
cosLookup[4421] <= 0.911498341;
cosLookup[4422] <= 0.911458901;
cosLookup[4423] <= 0.911419453;
cosLookup[4424] <= 0.911379996;
cosLookup[4425] <= 0.911340531;
cosLookup[4426] <= 0.911301058;
cosLookup[4427] <= 0.911261576;
cosLookup[4428] <= 0.911222086;
cosLookup[4429] <= 0.911182588;
cosLookup[4430] <= 0.911143081;
cosLookup[4431] <= 0.911103565;
cosLookup[4432] <= 0.911064042;
cosLookup[4433] <= 0.91102451;
cosLookup[4434] <= 0.910984969;
cosLookup[4435] <= 0.910945421;
cosLookup[4436] <= 0.910905864;
cosLookup[4437] <= 0.910866298;
cosLookup[4438] <= 0.910826724;
cosLookup[4439] <= 0.910787142;
cosLookup[4440] <= 0.910747551;
cosLookup[4441] <= 0.910707952;
cosLookup[4442] <= 0.910668345;
cosLookup[4443] <= 0.910628729;
cosLookup[4444] <= 0.910589105;
cosLookup[4445] <= 0.910549473;
cosLookup[4446] <= 0.910509832;
cosLookup[4447] <= 0.910470183;
cosLookup[4448] <= 0.910430525;
cosLookup[4449] <= 0.910390859;
cosLookup[4450] <= 0.910351185;
cosLookup[4451] <= 0.910311502;
cosLookup[4452] <= 0.910271811;
cosLookup[4453] <= 0.910232112;
cosLookup[4454] <= 0.910192404;
cosLookup[4455] <= 0.910152688;
cosLookup[4456] <= 0.910112963;
cosLookup[4457] <= 0.91007323;
cosLookup[4458] <= 0.910033489;
cosLookup[4459] <= 0.909993739;
cosLookup[4460] <= 0.909953981;
cosLookup[4461] <= 0.909914215;
cosLookup[4462] <= 0.90987444;
cosLookup[4463] <= 0.909834657;
cosLookup[4464] <= 0.909794866;
cosLookup[4465] <= 0.909755066;
cosLookup[4466] <= 0.909715258;
cosLookup[4467] <= 0.909675441;
cosLookup[4468] <= 0.909635616;
cosLookup[4469] <= 0.909595783;
cosLookup[4470] <= 0.909555941;
cosLookup[4471] <= 0.909516091;
cosLookup[4472] <= 0.909476233;
cosLookup[4473] <= 0.909436366;
cosLookup[4474] <= 0.909396491;
cosLookup[4475] <= 0.909356608;
cosLookup[4476] <= 0.909316716;
cosLookup[4477] <= 0.909276816;
cosLookup[4478] <= 0.909236907;
cosLookup[4479] <= 0.90919699;
cosLookup[4480] <= 0.909157065;
cosLookup[4481] <= 0.909117132;
cosLookup[4482] <= 0.90907719;
cosLookup[4483] <= 0.909037239;
cosLookup[4484] <= 0.908997281;
cosLookup[4485] <= 0.908957314;
cosLookup[4486] <= 0.908917338;
cosLookup[4487] <= 0.908877355;
cosLookup[4488] <= 0.908837363;
cosLookup[4489] <= 0.908797362;
cosLookup[4490] <= 0.908757353;
cosLookup[4491] <= 0.908717336;
cosLookup[4492] <= 0.908677311;
cosLookup[4493] <= 0.908637277;
cosLookup[4494] <= 0.908597235;
cosLookup[4495] <= 0.908557184;
cosLookup[4496] <= 0.908517125;
cosLookup[4497] <= 0.908477058;
cosLookup[4498] <= 0.908436982;
cosLookup[4499] <= 0.908396898;
cosLookup[4500] <= 0.908356806;
cosLookup[4501] <= 0.908316705;
cosLookup[4502] <= 0.908276596;
cosLookup[4503] <= 0.908236479;
cosLookup[4504] <= 0.908196353;
cosLookup[4505] <= 0.908156219;
cosLookup[4506] <= 0.908116077;
cosLookup[4507] <= 0.908075926;
cosLookup[4508] <= 0.908035767;
cosLookup[4509] <= 0.907995599;
cosLookup[4510] <= 0.907955424;
cosLookup[4511] <= 0.90791524;
cosLookup[4512] <= 0.907875047;
cosLookup[4513] <= 0.907834846;
cosLookup[4514] <= 0.907794637;
cosLookup[4515] <= 0.907754419;
cosLookup[4516] <= 0.907714194;
cosLookup[4517] <= 0.907673959;
cosLookup[4518] <= 0.907633717;
cosLookup[4519] <= 0.907593466;
cosLookup[4520] <= 0.907553207;
cosLookup[4521] <= 0.907512939;
cosLookup[4522] <= 0.907472663;
cosLookup[4523] <= 0.907432379;
cosLookup[4524] <= 0.907392086;
cosLookup[4525] <= 0.907351785;
cosLookup[4526] <= 0.907311476;
cosLookup[4527] <= 0.907271158;
cosLookup[4528] <= 0.907230832;
cosLookup[4529] <= 0.907190498;
cosLookup[4530] <= 0.907150155;
cosLookup[4531] <= 0.907109804;
cosLookup[4532] <= 0.907069445;
cosLookup[4533] <= 0.907029077;
cosLookup[4534] <= 0.906988701;
cosLookup[4535] <= 0.906948317;
cosLookup[4536] <= 0.906907924;
cosLookup[4537] <= 0.906867523;
cosLookup[4538] <= 0.906827114;
cosLookup[4539] <= 0.906786696;
cosLookup[4540] <= 0.90674627;
cosLookup[4541] <= 0.906705836;
cosLookup[4542] <= 0.906665393;
cosLookup[4543] <= 0.906624942;
cosLookup[4544] <= 0.906584483;
cosLookup[4545] <= 0.906544015;
cosLookup[4546] <= 0.906503539;
cosLookup[4547] <= 0.906463054;
cosLookup[4548] <= 0.906422562;
cosLookup[4549] <= 0.906382061;
cosLookup[4550] <= 0.906341551;
cosLookup[4551] <= 0.906301034;
cosLookup[4552] <= 0.906260507;
cosLookup[4553] <= 0.906219973;
cosLookup[4554] <= 0.90617943;
cosLookup[4555] <= 0.906138879;
cosLookup[4556] <= 0.90609832;
cosLookup[4557] <= 0.906057752;
cosLookup[4558] <= 0.906017176;
cosLookup[4559] <= 0.905976592;
cosLookup[4560] <= 0.905935999;
cosLookup[4561] <= 0.905895398;
cosLookup[4562] <= 0.905854789;
cosLookup[4563] <= 0.905814171;
cosLookup[4564] <= 0.905773545;
cosLookup[4565] <= 0.905732911;
cosLookup[4566] <= 0.905692268;
cosLookup[4567] <= 0.905651617;
cosLookup[4568] <= 0.905610958;
cosLookup[4569] <= 0.90557029;
cosLookup[4570] <= 0.905529614;
cosLookup[4571] <= 0.90548893;
cosLookup[4572] <= 0.905448237;
cosLookup[4573] <= 0.905407537;
cosLookup[4574] <= 0.905366827;
cosLookup[4575] <= 0.90532611;
cosLookup[4576] <= 0.905285384;
cosLookup[4577] <= 0.90524465;
cosLookup[4578] <= 0.905203907;
cosLookup[4579] <= 0.905163156;
cosLookup[4580] <= 0.905122397;
cosLookup[4581] <= 0.90508163;
cosLookup[4582] <= 0.905040854;
cosLookup[4583] <= 0.90500007;
cosLookup[4584] <= 0.904959277;
cosLookup[4585] <= 0.904918476;
cosLookup[4586] <= 0.904877667;
cosLookup[4587] <= 0.90483685;
cosLookup[4588] <= 0.904796024;
cosLookup[4589] <= 0.90475519;
cosLookup[4590] <= 0.904714348;
cosLookup[4591] <= 0.904673497;
cosLookup[4592] <= 0.904632638;
cosLookup[4593] <= 0.904591771;
cosLookup[4594] <= 0.904550895;
cosLookup[4595] <= 0.904510011;
cosLookup[4596] <= 0.904469119;
cosLookup[4597] <= 0.904428218;
cosLookup[4598] <= 0.904387309;
cosLookup[4599] <= 0.904346392;
cosLookup[4600] <= 0.904305467;
cosLookup[4601] <= 0.904264533;
cosLookup[4602] <= 0.904223591;
cosLookup[4603] <= 0.90418264;
cosLookup[4604] <= 0.904141681;
cosLookup[4605] <= 0.904100714;
cosLookup[4606] <= 0.904059739;
cosLookup[4607] <= 0.904018755;
cosLookup[4608] <= 0.903977763;
cosLookup[4609] <= 0.903936763;
cosLookup[4610] <= 0.903895754;
cosLookup[4611] <= 0.903854737;
cosLookup[4612] <= 0.903813712;
cosLookup[4613] <= 0.903772679;
cosLookup[4614] <= 0.903731637;
cosLookup[4615] <= 0.903690587;
cosLookup[4616] <= 0.903649528;
cosLookup[4617] <= 0.903608461;
cosLookup[4618] <= 0.903567386;
cosLookup[4619] <= 0.903526303;
cosLookup[4620] <= 0.903485211;
cosLookup[4621] <= 0.903444111;
cosLookup[4622] <= 0.903403003;
cosLookup[4623] <= 0.903361886;
cosLookup[4624] <= 0.903320761;
cosLookup[4625] <= 0.903279628;
cosLookup[4626] <= 0.903238486;
cosLookup[4627] <= 0.903197336;
cosLookup[4628] <= 0.903156178;
cosLookup[4629] <= 0.903115012;
cosLookup[4630] <= 0.903073837;
cosLookup[4631] <= 0.903032654;
cosLookup[4632] <= 0.902991463;
cosLookup[4633] <= 0.902950263;
cosLookup[4634] <= 0.902909055;
cosLookup[4635] <= 0.902867839;
cosLookup[4636] <= 0.902826614;
cosLookup[4637] <= 0.902785381;
cosLookup[4638] <= 0.90274414;
cosLookup[4639] <= 0.902702891;
cosLookup[4640] <= 0.902661633;
cosLookup[4641] <= 0.902620367;
cosLookup[4642] <= 0.902579093;
cosLookup[4643] <= 0.90253781;
cosLookup[4644] <= 0.902496519;
cosLookup[4645] <= 0.90245522;
cosLookup[4646] <= 0.902413912;
cosLookup[4647] <= 0.902372596;
cosLookup[4648] <= 0.902331272;
cosLookup[4649] <= 0.90228994;
cosLookup[4650] <= 0.902248599;
cosLookup[4651] <= 0.90220725;
cosLookup[4652] <= 0.902165893;
cosLookup[4653] <= 0.902124527;
cosLookup[4654] <= 0.902083153;
cosLookup[4655] <= 0.902041771;
cosLookup[4656] <= 0.902000381;
cosLookup[4657] <= 0.901958982;
cosLookup[4658] <= 0.901917575;
cosLookup[4659] <= 0.90187616;
cosLookup[4660] <= 0.901834736;
cosLookup[4661] <= 0.901793304;
cosLookup[4662] <= 0.901751864;
cosLookup[4663] <= 0.901710415;
cosLookup[4664] <= 0.901668958;
cosLookup[4665] <= 0.901627493;
cosLookup[4666] <= 0.90158602;
cosLookup[4667] <= 0.901544538;
cosLookup[4668] <= 0.901503048;
cosLookup[4669] <= 0.90146155;
cosLookup[4670] <= 0.901420044;
cosLookup[4671] <= 0.901378529;
cosLookup[4672] <= 0.901337006;
cosLookup[4673] <= 0.901295474;
cosLookup[4674] <= 0.901253935;
cosLookup[4675] <= 0.901212387;
cosLookup[4676] <= 0.90117083;
cosLookup[4677] <= 0.901129266;
cosLookup[4678] <= 0.901087693;
cosLookup[4679] <= 0.901046112;
cosLookup[4680] <= 0.901004523;
cosLookup[4681] <= 0.900962925;
cosLookup[4682] <= 0.900921319;
cosLookup[4683] <= 0.900879705;
cosLookup[4684] <= 0.900838082;
cosLookup[4685] <= 0.900796451;
cosLookup[4686] <= 0.900754812;
cosLookup[4687] <= 0.900713165;
cosLookup[4688] <= 0.900671509;
cosLookup[4689] <= 0.900629845;
cosLookup[4690] <= 0.900588173;
cosLookup[4691] <= 0.900546493;
cosLookup[4692] <= 0.900504804;
cosLookup[4693] <= 0.900463107;
cosLookup[4694] <= 0.900421402;
cosLookup[4695] <= 0.900379688;
cosLookup[4696] <= 0.900337966;
cosLookup[4697] <= 0.900296236;
cosLookup[4698] <= 0.900254498;
cosLookup[4699] <= 0.900212751;
cosLookup[4700] <= 0.900170996;
cosLookup[4701] <= 0.900129233;
cosLookup[4702] <= 0.900087461;
cosLookup[4703] <= 0.900045681;
cosLookup[4704] <= 0.900003893;
cosLookup[4705] <= 0.899962097;
cosLookup[4706] <= 0.899920292;
cosLookup[4707] <= 0.89987848;
cosLookup[4708] <= 0.899836658;
cosLookup[4709] <= 0.899794829;
cosLookup[4710] <= 0.899752991;
cosLookup[4711] <= 0.899711145;
cosLookup[4712] <= 0.899669291;
cosLookup[4713] <= 0.899627429;
cosLookup[4714] <= 0.899585558;
cosLookup[4715] <= 0.899543679;
cosLookup[4716] <= 0.899501791;
cosLookup[4717] <= 0.899459896;
cosLookup[4718] <= 0.899417992;
cosLookup[4719] <= 0.89937608;
cosLookup[4720] <= 0.899334159;
cosLookup[4721] <= 0.899292231;
cosLookup[4722] <= 0.899250294;
cosLookup[4723] <= 0.899208349;
cosLookup[4724] <= 0.899166395;
cosLookup[4725] <= 0.899124433;
cosLookup[4726] <= 0.899082463;
cosLookup[4727] <= 0.899040485;
cosLookup[4728] <= 0.898998499;
cosLookup[4729] <= 0.898956504;
cosLookup[4730] <= 0.898914501;
cosLookup[4731] <= 0.89887249;
cosLookup[4732] <= 0.89883047;
cosLookup[4733] <= 0.898788442;
cosLookup[4734] <= 0.898746406;
cosLookup[4735] <= 0.898704362;
cosLookup[4736] <= 0.898662309;
cosLookup[4737] <= 0.898620248;
cosLookup[4738] <= 0.898578179;
cosLookup[4739] <= 0.898536102;
cosLookup[4740] <= 0.898494016;
cosLookup[4741] <= 0.898451922;
cosLookup[4742] <= 0.89840982;
cosLookup[4743] <= 0.898367709;
cosLookup[4744] <= 0.898325591;
cosLookup[4745] <= 0.898283464;
cosLookup[4746] <= 0.898241328;
cosLookup[4747] <= 0.898199185;
cosLookup[4748] <= 0.898157033;
cosLookup[4749] <= 0.898114873;
cosLookup[4750] <= 0.898072705;
cosLookup[4751] <= 0.898030528;
cosLookup[4752] <= 0.897988344;
cosLookup[4753] <= 0.897946151;
cosLookup[4754] <= 0.897903949;
cosLookup[4755] <= 0.89786174;
cosLookup[4756] <= 0.897819522;
cosLookup[4757] <= 0.897777296;
cosLookup[4758] <= 0.897735062;
cosLookup[4759] <= 0.897692819;
cosLookup[4760] <= 0.897650568;
cosLookup[4761] <= 0.897608309;
cosLookup[4762] <= 0.897566042;
cosLookup[4763] <= 0.897523767;
cosLookup[4764] <= 0.897481483;
cosLookup[4765] <= 0.897439191;
cosLookup[4766] <= 0.89739689;
cosLookup[4767] <= 0.897354582;
cosLookup[4768] <= 0.897312265;
cosLookup[4769] <= 0.89726994;
cosLookup[4770] <= 0.897227607;
cosLookup[4771] <= 0.897185265;
cosLookup[4772] <= 0.897142915;
cosLookup[4773] <= 0.897100557;
cosLookup[4774] <= 0.897058191;
cosLookup[4775] <= 0.897015816;
cosLookup[4776] <= 0.896973434;
cosLookup[4777] <= 0.896931043;
cosLookup[4778] <= 0.896888643;
cosLookup[4779] <= 0.896846236;
cosLookup[4780] <= 0.89680382;
cosLookup[4781] <= 0.896761396;
cosLookup[4782] <= 0.896718964;
cosLookup[4783] <= 0.896676523;
cosLookup[4784] <= 0.896634075;
cosLookup[4785] <= 0.896591618;
cosLookup[4786] <= 0.896549152;
cosLookup[4787] <= 0.896506679;
cosLookup[4788] <= 0.896464197;
cosLookup[4789] <= 0.896421707;
cosLookup[4790] <= 0.896379209;
cosLookup[4791] <= 0.896336703;
cosLookup[4792] <= 0.896294188;
cosLookup[4793] <= 0.896251665;
cosLookup[4794] <= 0.896209134;
cosLookup[4795] <= 0.896166595;
cosLookup[4796] <= 0.896124047;
cosLookup[4797] <= 0.896081491;
cosLookup[4798] <= 0.896038927;
cosLookup[4799] <= 0.895996355;
cosLookup[4800] <= 0.895953774;
cosLookup[4801] <= 0.895911185;
cosLookup[4802] <= 0.895868588;
cosLookup[4803] <= 0.895825983;
cosLookup[4804] <= 0.895783369;
cosLookup[4805] <= 0.895740748;
cosLookup[4806] <= 0.895698118;
cosLookup[4807] <= 0.89565548;
cosLookup[4808] <= 0.895612833;
cosLookup[4809] <= 0.895570178;
cosLookup[4810] <= 0.895527515;
cosLookup[4811] <= 0.895484844;
cosLookup[4812] <= 0.895442165;
cosLookup[4813] <= 0.895399477;
cosLookup[4814] <= 0.895356781;
cosLookup[4815] <= 0.895314077;
cosLookup[4816] <= 0.895271365;
cosLookup[4817] <= 0.895228645;
cosLookup[4818] <= 0.895185916;
cosLookup[4819] <= 0.895143179;
cosLookup[4820] <= 0.895100434;
cosLookup[4821] <= 0.89505768;
cosLookup[4822] <= 0.895014918;
cosLookup[4823] <= 0.894972149;
cosLookup[4824] <= 0.89492937;
cosLookup[4825] <= 0.894886584;
cosLookup[4826] <= 0.894843789;
cosLookup[4827] <= 0.894800987;
cosLookup[4828] <= 0.894758176;
cosLookup[4829] <= 0.894715356;
cosLookup[4830] <= 0.894672529;
cosLookup[4831] <= 0.894629693;
cosLookup[4832] <= 0.894586849;
cosLookup[4833] <= 0.894543997;
cosLookup[4834] <= 0.894501137;
cosLookup[4835] <= 0.894458268;
cosLookup[4836] <= 0.894415391;
cosLookup[4837] <= 0.894372506;
cosLookup[4838] <= 0.894329613;
cosLookup[4839] <= 0.894286711;
cosLookup[4840] <= 0.894243802;
cosLookup[4841] <= 0.894200884;
cosLookup[4842] <= 0.894157957;
cosLookup[4843] <= 0.894115023;
cosLookup[4844] <= 0.894072081;
cosLookup[4845] <= 0.89402913;
cosLookup[4846] <= 0.893986171;
cosLookup[4847] <= 0.893943203;
cosLookup[4848] <= 0.893900228;
cosLookup[4849] <= 0.893857244;
cosLookup[4850] <= 0.893814252;
cosLookup[4851] <= 0.893771252;
cosLookup[4852] <= 0.893728244;
cosLookup[4853] <= 0.893685227;
cosLookup[4854] <= 0.893642203;
cosLookup[4855] <= 0.89359917;
cosLookup[4856] <= 0.893556128;
cosLookup[4857] <= 0.893513079;
cosLookup[4858] <= 0.893470021;
cosLookup[4859] <= 0.893426955;
cosLookup[4860] <= 0.893383881;
cosLookup[4861] <= 0.893340799;
cosLookup[4862] <= 0.893297709;
cosLookup[4863] <= 0.89325461;
cosLookup[4864] <= 0.893211503;
cosLookup[4865] <= 0.893168388;
cosLookup[4866] <= 0.893125265;
cosLookup[4867] <= 0.893082133;
cosLookup[4868] <= 0.893038993;
cosLookup[4869] <= 0.892995845;
cosLookup[4870] <= 0.892952689;
cosLookup[4871] <= 0.892909525;
cosLookup[4872] <= 0.892866352;
cosLookup[4873] <= 0.892823171;
cosLookup[4874] <= 0.892779982;
cosLookup[4875] <= 0.892736785;
cosLookup[4876] <= 0.89269358;
cosLookup[4877] <= 0.892650366;
cosLookup[4878] <= 0.892607144;
cosLookup[4879] <= 0.892563914;
cosLookup[4880] <= 0.892520676;
cosLookup[4881] <= 0.89247743;
cosLookup[4882] <= 0.892434175;
cosLookup[4883] <= 0.892390912;
cosLookup[4884] <= 0.892347641;
cosLookup[4885] <= 0.892304362;
cosLookup[4886] <= 0.892261074;
cosLookup[4887] <= 0.892217779;
cosLookup[4888] <= 0.892174475;
cosLookup[4889] <= 0.892131163;
cosLookup[4890] <= 0.892087842;
cosLookup[4891] <= 0.892044514;
cosLookup[4892] <= 0.892001177;
cosLookup[4893] <= 0.891957832;
cosLookup[4894] <= 0.891914479;
cosLookup[4895] <= 0.891871118;
cosLookup[4896] <= 0.891827749;
cosLookup[4897] <= 0.891784371;
cosLookup[4898] <= 0.891740985;
cosLookup[4899] <= 0.891697591;
cosLookup[4900] <= 0.891654189;
cosLookup[4901] <= 0.891610778;
cosLookup[4902] <= 0.89156736;
cosLookup[4903] <= 0.891523933;
cosLookup[4904] <= 0.891480498;
cosLookup[4905] <= 0.891437054;
cosLookup[4906] <= 0.891393603;
cosLookup[4907] <= 0.891350143;
cosLookup[4908] <= 0.891306675;
cosLookup[4909] <= 0.891263199;
cosLookup[4910] <= 0.891219715;
cosLookup[4911] <= 0.891176223;
cosLookup[4912] <= 0.891132722;
cosLookup[4913] <= 0.891089213;
cosLookup[4914] <= 0.891045696;
cosLookup[4915] <= 0.891002171;
cosLookup[4916] <= 0.890958638;
cosLookup[4917] <= 0.890915096;
cosLookup[4918] <= 0.890871547;
cosLookup[4919] <= 0.890827989;
cosLookup[4920] <= 0.890784423;
cosLookup[4921] <= 0.890740848;
cosLookup[4922] <= 0.890697266;
cosLookup[4923] <= 0.890653675;
cosLookup[4924] <= 0.890610076;
cosLookup[4925] <= 0.890566469;
cosLookup[4926] <= 0.890522854;
cosLookup[4927] <= 0.89047923;
cosLookup[4928] <= 0.890435599;
cosLookup[4929] <= 0.890391959;
cosLookup[4930] <= 0.890348311;
cosLookup[4931] <= 0.890304655;
cosLookup[4932] <= 0.89026099;
cosLookup[4933] <= 0.890217318;
cosLookup[4934] <= 0.890173637;
cosLookup[4935] <= 0.890129948;
cosLookup[4936] <= 0.890086251;
cosLookup[4937] <= 0.890042546;
cosLookup[4938] <= 0.889998832;
cosLookup[4939] <= 0.889955111;
cosLookup[4940] <= 0.889911381;
cosLookup[4941] <= 0.889867643;
cosLookup[4942] <= 0.889823897;
cosLookup[4943] <= 0.889780142;
cosLookup[4944] <= 0.88973638;
cosLookup[4945] <= 0.889692609;
cosLookup[4946] <= 0.88964883;
cosLookup[4947] <= 0.889605043;
cosLookup[4948] <= 0.889561248;
cosLookup[4949] <= 0.889517444;
cosLookup[4950] <= 0.889473633;
cosLookup[4951] <= 0.889429813;
cosLookup[4952] <= 0.889385985;
cosLookup[4953] <= 0.889342149;
cosLookup[4954] <= 0.889298305;
cosLookup[4955] <= 0.889254452;
cosLookup[4956] <= 0.889210591;
cosLookup[4957] <= 0.889166723;
cosLookup[4958] <= 0.889122846;
cosLookup[4959] <= 0.88907896;
cosLookup[4960] <= 0.889035067;
cosLookup[4961] <= 0.888991165;
cosLookup[4962] <= 0.888947256;
cosLookup[4963] <= 0.888903338;
cosLookup[4964] <= 0.888859412;
cosLookup[4965] <= 0.888815478;
cosLookup[4966] <= 0.888771535;
cosLookup[4967] <= 0.888727585;
cosLookup[4968] <= 0.888683626;
cosLookup[4969] <= 0.888639659;
cosLookup[4970] <= 0.888595684;
cosLookup[4971] <= 0.888551701;
cosLookup[4972] <= 0.888507709;
cosLookup[4973] <= 0.88846371;
cosLookup[4974] <= 0.888419702;
cosLookup[4975] <= 0.888375686;
cosLookup[4976] <= 0.888331662;
cosLookup[4977] <= 0.88828763;
cosLookup[4978] <= 0.888243589;
cosLookup[4979] <= 0.888199541;
cosLookup[4980] <= 0.888155484;
cosLookup[4981] <= 0.888111419;
cosLookup[4982] <= 0.888067346;
cosLookup[4983] <= 0.888023265;
cosLookup[4984] <= 0.887979175;
cosLookup[4985] <= 0.887935078;
cosLookup[4986] <= 0.887890972;
cosLookup[4987] <= 0.887846858;
cosLookup[4988] <= 0.887802736;
cosLookup[4989] <= 0.887758606;
cosLookup[4990] <= 0.887714467;
cosLookup[4991] <= 0.887670321;
cosLookup[4992] <= 0.887626166;
cosLookup[4993] <= 0.887582003;
cosLookup[4994] <= 0.887537832;
cosLookup[4995] <= 0.887493653;
cosLookup[4996] <= 0.887449466;
cosLookup[4997] <= 0.88740527;
cosLookup[4998] <= 0.887361067;
cosLookup[4999] <= 0.887316855;
cosLookup[5000] <= 0.887272635;
cosLookup[5001] <= 0.887228407;
cosLookup[5002] <= 0.88718417;
cosLookup[5003] <= 0.887139926;
cosLookup[5004] <= 0.887095673;
cosLookup[5005] <= 0.887051413;
cosLookup[5006] <= 0.887007144;
cosLookup[5007] <= 0.886962867;
cosLookup[5008] <= 0.886918582;
cosLookup[5009] <= 0.886874288;
cosLookup[5010] <= 0.886829987;
cosLookup[5011] <= 0.886785677;
cosLookup[5012] <= 0.886741359;
cosLookup[5013] <= 0.886697033;
cosLookup[5014] <= 0.886652699;
cosLookup[5015] <= 0.886608357;
cosLookup[5016] <= 0.886564006;
cosLookup[5017] <= 0.886519648;
cosLookup[5018] <= 0.886475281;
cosLookup[5019] <= 0.886430906;
cosLookup[5020] <= 0.886386523;
cosLookup[5021] <= 0.886342132;
cosLookup[5022] <= 0.886297733;
cosLookup[5023] <= 0.886253325;
cosLookup[5024] <= 0.88620891;
cosLookup[5025] <= 0.886164486;
cosLookup[5026] <= 0.886120054;
cosLookup[5027] <= 0.886075614;
cosLookup[5028] <= 0.886031166;
cosLookup[5029] <= 0.885986709;
cosLookup[5030] <= 0.885942245;
cosLookup[5031] <= 0.885897772;
cosLookup[5032] <= 0.885853292;
cosLookup[5033] <= 0.885808803;
cosLookup[5034] <= 0.885764306;
cosLookup[5035] <= 0.8857198;
cosLookup[5036] <= 0.885675287;
cosLookup[5037] <= 0.885630765;
cosLookup[5038] <= 0.885586236;
cosLookup[5039] <= 0.885541698;
cosLookup[5040] <= 0.885497152;
cosLookup[5041] <= 0.885452598;
cosLookup[5042] <= 0.885408036;
cosLookup[5043] <= 0.885363466;
cosLookup[5044] <= 0.885318887;
cosLookup[5045] <= 0.885274301;
cosLookup[5046] <= 0.885229706;
cosLookup[5047] <= 0.885185103;
cosLookup[5048] <= 0.885140492;
cosLookup[5049] <= 0.885095873;
cosLookup[5050] <= 0.885051245;
cosLookup[5051] <= 0.88500661;
cosLookup[5052] <= 0.884961966;
cosLookup[5053] <= 0.884917315;
cosLookup[5054] <= 0.884872655;
cosLookup[5055] <= 0.884827987;
cosLookup[5056] <= 0.884783311;
cosLookup[5057] <= 0.884738627;
cosLookup[5058] <= 0.884693934;
cosLookup[5059] <= 0.884649234;
cosLookup[5060] <= 0.884604525;
cosLookup[5061] <= 0.884559808;
cosLookup[5062] <= 0.884515083;
cosLookup[5063] <= 0.88447035;
cosLookup[5064] <= 0.884425609;
cosLookup[5065] <= 0.88438086;
cosLookup[5066] <= 0.884336102;
cosLookup[5067] <= 0.884291337;
cosLookup[5068] <= 0.884246563;
cosLookup[5069] <= 0.884201781;
cosLookup[5070] <= 0.884156991;
cosLookup[5071] <= 0.884112193;
cosLookup[5072] <= 0.884067387;
cosLookup[5073] <= 0.884022573;
cosLookup[5074] <= 0.88397775;
cosLookup[5075] <= 0.88393292;
cosLookup[5076] <= 0.883888081;
cosLookup[5077] <= 0.883843234;
cosLookup[5078] <= 0.883798379;
cosLookup[5079] <= 0.883753516;
cosLookup[5080] <= 0.883708645;
cosLookup[5081] <= 0.883663766;
cosLookup[5082] <= 0.883618878;
cosLookup[5083] <= 0.883573983;
cosLookup[5084] <= 0.883529079;
cosLookup[5085] <= 0.883484167;
cosLookup[5086] <= 0.883439247;
cosLookup[5087] <= 0.883394319;
cosLookup[5088] <= 0.883349383;
cosLookup[5089] <= 0.883304439;
cosLookup[5090] <= 0.883259486;
cosLookup[5091] <= 0.883214526;
cosLookup[5092] <= 0.883169557;
cosLookup[5093] <= 0.88312458;
cosLookup[5094] <= 0.883079595;
cosLookup[5095] <= 0.883034602;
cosLookup[5096] <= 0.882989601;
cosLookup[5097] <= 0.882944592;
cosLookup[5098] <= 0.882899575;
cosLookup[5099] <= 0.882854549;
cosLookup[5100] <= 0.882809516;
cosLookup[5101] <= 0.882764474;
cosLookup[5102] <= 0.882719424;
cosLookup[5103] <= 0.882674366;
cosLookup[5104] <= 0.8826293;
cosLookup[5105] <= 0.882584226;
cosLookup[5106] <= 0.882539144;
cosLookup[5107] <= 0.882494053;
cosLookup[5108] <= 0.882448955;
cosLookup[5109] <= 0.882403848;
cosLookup[5110] <= 0.882358733;
cosLookup[5111] <= 0.88231361;
cosLookup[5112] <= 0.882268479;
cosLookup[5113] <= 0.88222334;
cosLookup[5114] <= 0.882178193;
cosLookup[5115] <= 0.882133038;
cosLookup[5116] <= 0.882087874;
cosLookup[5117] <= 0.882042703;
cosLookup[5118] <= 0.881997523;
cosLookup[5119] <= 0.881952336;
cosLookup[5120] <= 0.88190714;
cosLookup[5121] <= 0.881861936;
cosLookup[5122] <= 0.881816724;
cosLookup[5123] <= 0.881771504;
cosLookup[5124] <= 0.881726275;
cosLookup[5125] <= 0.881681039;
cosLookup[5126] <= 0.881635795;
cosLookup[5127] <= 0.881590542;
cosLookup[5128] <= 0.881545281;
cosLookup[5129] <= 0.881500012;
cosLookup[5130] <= 0.881454736;
cosLookup[5131] <= 0.881409451;
cosLookup[5132] <= 0.881364158;
cosLookup[5133] <= 0.881318856;
cosLookup[5134] <= 0.881273547;
cosLookup[5135] <= 0.88122823;
cosLookup[5136] <= 0.881182904;
cosLookup[5137] <= 0.881137571;
cosLookup[5138] <= 0.881092229;
cosLookup[5139] <= 0.881046879;
cosLookup[5140] <= 0.881001521;
cosLookup[5141] <= 0.880956155;
cosLookup[5142] <= 0.880910781;
cosLookup[5143] <= 0.880865399;
cosLookup[5144] <= 0.880820009;
cosLookup[5145] <= 0.88077461;
cosLookup[5146] <= 0.880729204;
cosLookup[5147] <= 0.880683789;
cosLookup[5148] <= 0.880638366;
cosLookup[5149] <= 0.880592936;
cosLookup[5150] <= 0.880547497;
cosLookup[5151] <= 0.88050205;
cosLookup[5152] <= 0.880456595;
cosLookup[5153] <= 0.880411132;
cosLookup[5154] <= 0.88036566;
cosLookup[5155] <= 0.880320181;
cosLookup[5156] <= 0.880274694;
cosLookup[5157] <= 0.880229198;
cosLookup[5158] <= 0.880183694;
cosLookup[5159] <= 0.880138183;
cosLookup[5160] <= 0.880092663;
cosLookup[5161] <= 0.880047135;
cosLookup[5162] <= 0.880001599;
cosLookup[5163] <= 0.879956055;
cosLookup[5164] <= 0.879910503;
cosLookup[5165] <= 0.879864942;
cosLookup[5166] <= 0.879819374;
cosLookup[5167] <= 0.879773798;
cosLookup[5168] <= 0.879728213;
cosLookup[5169] <= 0.879682621;
cosLookup[5170] <= 0.87963702;
cosLookup[5171] <= 0.879591411;
cosLookup[5172] <= 0.879545794;
cosLookup[5173] <= 0.879500169;
cosLookup[5174] <= 0.879454536;
cosLookup[5175] <= 0.879408895;
cosLookup[5176] <= 0.879363246;
cosLookup[5177] <= 0.879317589;
cosLookup[5178] <= 0.879271923;
cosLookup[5179] <= 0.87922625;
cosLookup[5180] <= 0.879180568;
cosLookup[5181] <= 0.879134879;
cosLookup[5182] <= 0.879089181;
cosLookup[5183] <= 0.879043475;
cosLookup[5184] <= 0.878997761;
cosLookup[5185] <= 0.878952039;
cosLookup[5186] <= 0.878906309;
cosLookup[5187] <= 0.878860571;
cosLookup[5188] <= 0.878814825;
cosLookup[5189] <= 0.878769071;
cosLookup[5190] <= 0.878723309;
cosLookup[5191] <= 0.878677538;
cosLookup[5192] <= 0.87863176;
cosLookup[5193] <= 0.878585973;
cosLookup[5194] <= 0.878540178;
cosLookup[5195] <= 0.878494376;
cosLookup[5196] <= 0.878448565;
cosLookup[5197] <= 0.878402746;
cosLookup[5198] <= 0.878356919;
cosLookup[5199] <= 0.878311084;
cosLookup[5200] <= 0.878265241;
cosLookup[5201] <= 0.87821939;
cosLookup[5202] <= 0.878173531;
cosLookup[5203] <= 0.878127663;
cosLookup[5204] <= 0.878081788;
cosLookup[5205] <= 0.878035904;
cosLookup[5206] <= 0.877990013;
cosLookup[5207] <= 0.877944113;
cosLookup[5208] <= 0.877898206;
cosLookup[5209] <= 0.87785229;
cosLookup[5210] <= 0.877806366;
cosLookup[5211] <= 0.877760434;
cosLookup[5212] <= 0.877714494;
cosLookup[5213] <= 0.877668546;
cosLookup[5214] <= 0.87762259;
cosLookup[5215] <= 0.877576626;
cosLookup[5216] <= 0.877530654;
cosLookup[5217] <= 0.877484673;
cosLookup[5218] <= 0.877438685;
cosLookup[5219] <= 0.877392689;
cosLookup[5220] <= 0.877346684;
cosLookup[5221] <= 0.877300671;
cosLookup[5222] <= 0.877254651;
cosLookup[5223] <= 0.877208622;
cosLookup[5224] <= 0.877162585;
cosLookup[5225] <= 0.877116541;
cosLookup[5226] <= 0.877070488;
cosLookup[5227] <= 0.877024427;
cosLookup[5228] <= 0.876978358;
cosLookup[5229] <= 0.876932281;
cosLookup[5230] <= 0.876886196;
cosLookup[5231] <= 0.876840102;
cosLookup[5232] <= 0.876794001;
cosLookup[5233] <= 0.876747892;
cosLookup[5234] <= 0.876701774;
cosLookup[5235] <= 0.876655649;
cosLookup[5236] <= 0.876609516;
cosLookup[5237] <= 0.876563374;
cosLookup[5238] <= 0.876517224;
cosLookup[5239] <= 0.876471067;
cosLookup[5240] <= 0.876424901;
cosLookup[5241] <= 0.876378727;
cosLookup[5242] <= 0.876332545;
cosLookup[5243] <= 0.876286355;
cosLookup[5244] <= 0.876240158;
cosLookup[5245] <= 0.876193952;
cosLookup[5246] <= 0.876147737;
cosLookup[5247] <= 0.876101515;
cosLookup[5248] <= 0.876055285;
cosLookup[5249] <= 0.876009047;
cosLookup[5250] <= 0.875962801;
cosLookup[5251] <= 0.875916546;
cosLookup[5252] <= 0.875870284;
cosLookup[5253] <= 0.875824014;
cosLookup[5254] <= 0.875777735;
cosLookup[5255] <= 0.875731449;
cosLookup[5256] <= 0.875685154;
cosLookup[5257] <= 0.875638851;
cosLookup[5258] <= 0.875592541;
cosLookup[5259] <= 0.875546222;
cosLookup[5260] <= 0.875499895;
cosLookup[5261] <= 0.87545356;
cosLookup[5262] <= 0.875407217;
cosLookup[5263] <= 0.875360867;
cosLookup[5264] <= 0.875314508;
cosLookup[5265] <= 0.875268141;
cosLookup[5266] <= 0.875221766;
cosLookup[5267] <= 0.875175382;
cosLookup[5268] <= 0.875128991;
cosLookup[5269] <= 0.875082592;
cosLookup[5270] <= 0.875036185;
cosLookup[5271] <= 0.87498977;
cosLookup[5272] <= 0.874943346;
cosLookup[5273] <= 0.874896915;
cosLookup[5274] <= 0.874850475;
cosLookup[5275] <= 0.874804028;
cosLookup[5276] <= 0.874757572;
cosLookup[5277] <= 0.874711109;
cosLookup[5278] <= 0.874664637;
cosLookup[5279] <= 0.874618158;
cosLookup[5280] <= 0.87457167;
cosLookup[5281] <= 0.874525174;
cosLookup[5282] <= 0.874478671;
cosLookup[5283] <= 0.874432159;
cosLookup[5284] <= 0.874385639;
cosLookup[5285] <= 0.874339111;
cosLookup[5286] <= 0.874292575;
cosLookup[5287] <= 0.874246031;
cosLookup[5288] <= 0.874199479;
cosLookup[5289] <= 0.874152919;
cosLookup[5290] <= 0.874106351;
cosLookup[5291] <= 0.874059775;
cosLookup[5292] <= 0.874013191;
cosLookup[5293] <= 0.873966599;
cosLookup[5294] <= 0.873919999;
cosLookup[5295] <= 0.87387339;
cosLookup[5296] <= 0.873826774;
cosLookup[5297] <= 0.87378015;
cosLookup[5298] <= 0.873733518;
cosLookup[5299] <= 0.873686877;
cosLookup[5300] <= 0.873640229;
cosLookup[5301] <= 0.873593573;
cosLookup[5302] <= 0.873546908;
cosLookup[5303] <= 0.873500236;
cosLookup[5304] <= 0.873453555;
cosLookup[5305] <= 0.873406867;
cosLookup[5306] <= 0.87336017;
cosLookup[5307] <= 0.873313465;
cosLookup[5308] <= 0.873266753;
cosLookup[5309] <= 0.873220032;
cosLookup[5310] <= 0.873173303;
cosLookup[5311] <= 0.873126567;
cosLookup[5312] <= 0.873079822;
cosLookup[5313] <= 0.873033069;
cosLookup[5314] <= 0.872986308;
cosLookup[5315] <= 0.87293954;
cosLookup[5316] <= 0.872892763;
cosLookup[5317] <= 0.872845978;
cosLookup[5318] <= 0.872799185;
cosLookup[5319] <= 0.872752384;
cosLookup[5320] <= 0.872705575;
cosLookup[5321] <= 0.872658758;
cosLookup[5322] <= 0.872611933;
cosLookup[5323] <= 0.8725651;
cosLookup[5324] <= 0.872518259;
cosLookup[5325] <= 0.87247141;
cosLookup[5326] <= 0.872424553;
cosLookup[5327] <= 0.872377688;
cosLookup[5328] <= 0.872330815;
cosLookup[5329] <= 0.872283934;
cosLookup[5330] <= 0.872237045;
cosLookup[5331] <= 0.872190148;
cosLookup[5332] <= 0.872143243;
cosLookup[5333] <= 0.872096329;
cosLookup[5334] <= 0.872049408;
cosLookup[5335] <= 0.872002479;
cosLookup[5336] <= 0.871955542;
cosLookup[5337] <= 0.871908596;
cosLookup[5338] <= 0.871861643;
cosLookup[5339] <= 0.871814682;
cosLookup[5340] <= 0.871767713;
cosLookup[5341] <= 0.871720735;
cosLookup[5342] <= 0.87167375;
cosLookup[5343] <= 0.871626757;
cosLookup[5344] <= 0.871579755;
cosLookup[5345] <= 0.871532746;
cosLookup[5346] <= 0.871485729;
cosLookup[5347] <= 0.871438703;
cosLookup[5348] <= 0.87139167;
cosLookup[5349] <= 0.871344628;
cosLookup[5350] <= 0.871297579;
cosLookup[5351] <= 0.871250521;
cosLookup[5352] <= 0.871203456;
cosLookup[5353] <= 0.871156383;
cosLookup[5354] <= 0.871109301;
cosLookup[5355] <= 0.871062212;
cosLookup[5356] <= 0.871015114;
cosLookup[5357] <= 0.870968009;
cosLookup[5358] <= 0.870920895;
cosLookup[5359] <= 0.870873774;
cosLookup[5360] <= 0.870826644;
cosLookup[5361] <= 0.870779507;
cosLookup[5362] <= 0.870732361;
cosLookup[5363] <= 0.870685208;
cosLookup[5364] <= 0.870638046;
cosLookup[5365] <= 0.870590877;
cosLookup[5366] <= 0.870543699;
cosLookup[5367] <= 0.870496514;
cosLookup[5368] <= 0.87044932;
cosLookup[5369] <= 0.870402119;
cosLookup[5370] <= 0.870354909;
cosLookup[5371] <= 0.870307692;
cosLookup[5372] <= 0.870260466;
cosLookup[5373] <= 0.870213232;
cosLookup[5374] <= 0.870165991;
cosLookup[5375] <= 0.870118741;
cosLookup[5376] <= 0.870071484;
cosLookup[5377] <= 0.870024218;
cosLookup[5378] <= 0.869976945;
cosLookup[5379] <= 0.869929663;
cosLookup[5380] <= 0.869882374;
cosLookup[5381] <= 0.869835076;
cosLookup[5382] <= 0.869787771;
cosLookup[5383] <= 0.869740457;
cosLookup[5384] <= 0.869693136;
cosLookup[5385] <= 0.869645806;
cosLookup[5386] <= 0.869598469;
cosLookup[5387] <= 0.869551123;
cosLookup[5388] <= 0.86950377;
cosLookup[5389] <= 0.869456408;
cosLookup[5390] <= 0.869409039;
cosLookup[5391] <= 0.869361661;
cosLookup[5392] <= 0.869314276;
cosLookup[5393] <= 0.869266882;
cosLookup[5394] <= 0.869219481;
cosLookup[5395] <= 0.869172072;
cosLookup[5396] <= 0.869124654;
cosLookup[5397] <= 0.869077229;
cosLookup[5398] <= 0.869029795;
cosLookup[5399] <= 0.868982354;
cosLookup[5400] <= 0.868934905;
cosLookup[5401] <= 0.868887447;
cosLookup[5402] <= 0.868839982;
cosLookup[5403] <= 0.868792508;
cosLookup[5404] <= 0.868745027;
cosLookup[5405] <= 0.868697538;
cosLookup[5406] <= 0.868650041;
cosLookup[5407] <= 0.868602535;
cosLookup[5408] <= 0.868555022;
cosLookup[5409] <= 0.868507501;
cosLookup[5410] <= 0.868459972;
cosLookup[5411] <= 0.868412434;
cosLookup[5412] <= 0.868364889;
cosLookup[5413] <= 0.868317336;
cosLookup[5414] <= 0.868269775;
cosLookup[5415] <= 0.868222206;
cosLookup[5416] <= 0.868174628;
cosLookup[5417] <= 0.868127043;
cosLookup[5418] <= 0.86807945;
cosLookup[5419] <= 0.868031849;
cosLookup[5420] <= 0.86798424;
cosLookup[5421] <= 0.867936623;
cosLookup[5422] <= 0.867888998;
cosLookup[5423] <= 0.867841365;
cosLookup[5424] <= 0.867793724;
cosLookup[5425] <= 0.867746075;
cosLookup[5426] <= 0.867698418;
cosLookup[5427] <= 0.867650753;
cosLookup[5428] <= 0.86760308;
cosLookup[5429] <= 0.8675554;
cosLookup[5430] <= 0.867507711;
cosLookup[5431] <= 0.867460014;
cosLookup[5432] <= 0.867412309;
cosLookup[5433] <= 0.867364596;
cosLookup[5434] <= 0.867316876;
cosLookup[5435] <= 0.867269147;
cosLookup[5436] <= 0.86722141;
cosLookup[5437] <= 0.867173666;
cosLookup[5438] <= 0.867125913;
cosLookup[5439] <= 0.867078153;
cosLookup[5440] <= 0.867030384;
cosLookup[5441] <= 0.866982607;
cosLookup[5442] <= 0.866934823;
cosLookup[5443] <= 0.86688703;
cosLookup[5444] <= 0.86683923;
cosLookup[5445] <= 0.866791422;
cosLookup[5446] <= 0.866743605;
cosLookup[5447] <= 0.866695781;
cosLookup[5448] <= 0.866647949;
cosLookup[5449] <= 0.866600108;
cosLookup[5450] <= 0.86655226;
cosLookup[5451] <= 0.866504404;
cosLookup[5452] <= 0.86645654;
cosLookup[5453] <= 0.866408668;
cosLookup[5454] <= 0.866360787;
cosLookup[5455] <= 0.866312899;
cosLookup[5456] <= 0.866265003;
cosLookup[5457] <= 0.866217099;
cosLookup[5458] <= 0.866169187;
cosLookup[5459] <= 0.866121268;
cosLookup[5460] <= 0.86607334;
cosLookup[5461] <= 0.866025404;
cosLookup[5462] <= 0.86597746;
cosLookup[5463] <= 0.865929508;
cosLookup[5464] <= 0.865881548;
cosLookup[5465] <= 0.865833581;
cosLookup[5466] <= 0.865785605;
cosLookup[5467] <= 0.865737622;
cosLookup[5468] <= 0.86568963;
cosLookup[5469] <= 0.86564163;
cosLookup[5470] <= 0.865593623;
cosLookup[5471] <= 0.865545608;
cosLookup[5472] <= 0.865497584;
cosLookup[5473] <= 0.865449553;
cosLookup[5474] <= 0.865401513;
cosLookup[5475] <= 0.865353466;
cosLookup[5476] <= 0.865305411;
cosLookup[5477] <= 0.865257348;
cosLookup[5478] <= 0.865209277;
cosLookup[5479] <= 0.865161198;
cosLookup[5480] <= 0.865113111;
cosLookup[5481] <= 0.865065016;
cosLookup[5482] <= 0.865016913;
cosLookup[5483] <= 0.864968802;
cosLookup[5484] <= 0.864920683;
cosLookup[5485] <= 0.864872556;
cosLookup[5486] <= 0.864824421;
cosLookup[5487] <= 0.864776279;
cosLookup[5488] <= 0.864728128;
cosLookup[5489] <= 0.864679969;
cosLookup[5490] <= 0.864631803;
cosLookup[5491] <= 0.864583628;
cosLookup[5492] <= 0.864535446;
cosLookup[5493] <= 0.864487256;
cosLookup[5494] <= 0.864439057;
cosLookup[5495] <= 0.864390851;
cosLookup[5496] <= 0.864342637;
cosLookup[5497] <= 0.864294415;
cosLookup[5498] <= 0.864246184;
cosLookup[5499] <= 0.864197946;
cosLookup[5500] <= 0.8641497;
cosLookup[5501] <= 0.864101446;
cosLookup[5502] <= 0.864053185;
cosLookup[5503] <= 0.864004915;
cosLookup[5504] <= 0.863956637;
cosLookup[5505] <= 0.863908351;
cosLookup[5506] <= 0.863860058;
cosLookup[5507] <= 0.863811756;
cosLookup[5508] <= 0.863763446;
cosLookup[5509] <= 0.863715129;
cosLookup[5510] <= 0.863666803;
cosLookup[5511] <= 0.86361847;
cosLookup[5512] <= 0.863570129;
cosLookup[5513] <= 0.86352178;
cosLookup[5514] <= 0.863473422;
cosLookup[5515] <= 0.863425057;
cosLookup[5516] <= 0.863376684;
cosLookup[5517] <= 0.863328303;
cosLookup[5518] <= 0.863279914;
cosLookup[5519] <= 0.863231517;
cosLookup[5520] <= 0.863183113;
cosLookup[5521] <= 0.8631347;
cosLookup[5522] <= 0.863086279;
cosLookup[5523] <= 0.863037851;
cosLookup[5524] <= 0.862989414;
cosLookup[5525] <= 0.86294097;
cosLookup[5526] <= 0.862892517;
cosLookup[5527] <= 0.862844057;
cosLookup[5528] <= 0.862795589;
cosLookup[5529] <= 0.862747112;
cosLookup[5530] <= 0.862698628;
cosLookup[5531] <= 0.862650136;
cosLookup[5532] <= 0.862601636;
cosLookup[5533] <= 0.862553128;
cosLookup[5534] <= 0.862504612;
cosLookup[5535] <= 0.862456089;
cosLookup[5536] <= 0.862407557;
cosLookup[5537] <= 0.862359017;
cosLookup[5538] <= 0.86231047;
cosLookup[5539] <= 0.862261914;
cosLookup[5540] <= 0.862213351;
cosLookup[5541] <= 0.862164779;
cosLookup[5542] <= 0.8621162;
cosLookup[5543] <= 0.862067613;
cosLookup[5544] <= 0.862019018;
cosLookup[5545] <= 0.861970415;
cosLookup[5546] <= 0.861921804;
cosLookup[5547] <= 0.861873185;
cosLookup[5548] <= 0.861824558;
cosLookup[5549] <= 0.861775923;
cosLookup[5550] <= 0.861727281;
cosLookup[5551] <= 0.86167863;
cosLookup[5552] <= 0.861629971;
cosLookup[5553] <= 0.861581305;
cosLookup[5554] <= 0.861532631;
cosLookup[5555] <= 0.861483948;
cosLookup[5556] <= 0.861435258;
cosLookup[5557] <= 0.86138656;
cosLookup[5558] <= 0.861337854;
cosLookup[5559] <= 0.86128914;
cosLookup[5560] <= 0.861240418;
cosLookup[5561] <= 0.861191689;
cosLookup[5562] <= 0.861142951;
cosLookup[5563] <= 0.861094205;
cosLookup[5564] <= 0.861045452;
cosLookup[5565] <= 0.86099669;
cosLookup[5566] <= 0.860947921;
cosLookup[5567] <= 0.860899144;
cosLookup[5568] <= 0.860850358;
cosLookup[5569] <= 0.860801565;
cosLookup[5570] <= 0.860752764;
cosLookup[5571] <= 0.860703955;
cosLookup[5572] <= 0.860655139;
cosLookup[5573] <= 0.860606314;
cosLookup[5574] <= 0.860557481;
cosLookup[5575] <= 0.860508641;
cosLookup[5576] <= 0.860459792;
cosLookup[5577] <= 0.860410936;
cosLookup[5578] <= 0.860362071;
cosLookup[5579] <= 0.860313199;
cosLookup[5580] <= 0.860264319;
cosLookup[5581] <= 0.860215431;
cosLookup[5582] <= 0.860166535;
cosLookup[5583] <= 0.860117631;
cosLookup[5584] <= 0.860068719;
cosLookup[5585] <= 0.8600198;
cosLookup[5586] <= 0.859970872;
cosLookup[5587] <= 0.859921937;
cosLookup[5588] <= 0.859872993;
cosLookup[5589] <= 0.859824042;
cosLookup[5590] <= 0.859775083;
cosLookup[5591] <= 0.859726116;
cosLookup[5592] <= 0.859677141;
cosLookup[5593] <= 0.859628158;
cosLookup[5594] <= 0.859579167;
cosLookup[5595] <= 0.859530168;
cosLookup[5596] <= 0.859481162;
cosLookup[5597] <= 0.859432147;
cosLookup[5598] <= 0.859383125;
cosLookup[5599] <= 0.859334095;
cosLookup[5600] <= 0.859285056;
cosLookup[5601] <= 0.85923601;
cosLookup[5602] <= 0.859186956;
cosLookup[5603] <= 0.859137894;
cosLookup[5604] <= 0.859088825;
cosLookup[5605] <= 0.859039747;
cosLookup[5606] <= 0.858990661;
cosLookup[5607] <= 0.858941568;
cosLookup[5608] <= 0.858892466;
cosLookup[5609] <= 0.858843357;
cosLookup[5610] <= 0.85879424;
cosLookup[5611] <= 0.858745115;
cosLookup[5612] <= 0.858695982;
cosLookup[5613] <= 0.858646841;
cosLookup[5614] <= 0.858597692;
cosLookup[5615] <= 0.858548536;
cosLookup[5616] <= 0.858499371;
cosLookup[5617] <= 0.858450199;
cosLookup[5618] <= 0.858401018;
cosLookup[5619] <= 0.85835183;
cosLookup[5620] <= 0.858302634;
cosLookup[5621] <= 0.85825343;
cosLookup[5622] <= 0.858204218;
cosLookup[5623] <= 0.858154998;
cosLookup[5624] <= 0.858105771;
cosLookup[5625] <= 0.858056535;
cosLookup[5626] <= 0.858007292;
cosLookup[5627] <= 0.85795804;
cosLookup[5628] <= 0.857908781;
cosLookup[5629] <= 0.857859514;
cosLookup[5630] <= 0.857810239;
cosLookup[5631] <= 0.857760956;
cosLookup[5632] <= 0.857711665;
cosLookup[5633] <= 0.857662367;
cosLookup[5634] <= 0.85761306;
cosLookup[5635] <= 0.857563746;
cosLookup[5636] <= 0.857514424;
cosLookup[5637] <= 0.857465093;
cosLookup[5638] <= 0.857415755;
cosLookup[5639] <= 0.857366409;
cosLookup[5640] <= 0.857317056;
cosLookup[5641] <= 0.857267694;
cosLookup[5642] <= 0.857218324;
cosLookup[5643] <= 0.857168947;
cosLookup[5644] <= 0.857119561;
cosLookup[5645] <= 0.857070168;
cosLookup[5646] <= 0.857020767;
cosLookup[5647] <= 0.856971358;
cosLookup[5648] <= 0.856921941;
cosLookup[5649] <= 0.856872516;
cosLookup[5650] <= 0.856823084;
cosLookup[5651] <= 0.856773643;
cosLookup[5652] <= 0.856724195;
cosLookup[5653] <= 0.856674739;
cosLookup[5654] <= 0.856625275;
cosLookup[5655] <= 0.856575803;
cosLookup[5656] <= 0.856526323;
cosLookup[5657] <= 0.856476835;
cosLookup[5658] <= 0.856427339;
cosLookup[5659] <= 0.856377836;
cosLookup[5660] <= 0.856328325;
cosLookup[5661] <= 0.856278805;
cosLookup[5662] <= 0.856229278;
cosLookup[5663] <= 0.856179743;
cosLookup[5664] <= 0.8561302;
cosLookup[5665] <= 0.85608065;
cosLookup[5666] <= 0.856031091;
cosLookup[5667] <= 0.855981525;
cosLookup[5668] <= 0.85593195;
cosLookup[5669] <= 0.855882368;
cosLookup[5670] <= 0.855832778;
cosLookup[5671] <= 0.85578318;
cosLookup[5672] <= 0.855733574;
cosLookup[5673] <= 0.855683961;
cosLookup[5674] <= 0.855634339;
cosLookup[5675] <= 0.85558471;
cosLookup[5676] <= 0.855535072;
cosLookup[5677] <= 0.855485427;
cosLookup[5678] <= 0.855435774;
cosLookup[5679] <= 0.855386113;
cosLookup[5680] <= 0.855336445;
cosLookup[5681] <= 0.855286768;
cosLookup[5682] <= 0.855237084;
cosLookup[5683] <= 0.855187391;
cosLookup[5684] <= 0.855137691;
cosLookup[5685] <= 0.855087983;
cosLookup[5686] <= 0.855038267;
cosLookup[5687] <= 0.854988544;
cosLookup[5688] <= 0.854938812;
cosLookup[5689] <= 0.854889072;
cosLookup[5690] <= 0.854839325;
cosLookup[5691] <= 0.85478957;
cosLookup[5692] <= 0.854739807;
cosLookup[5693] <= 0.854690036;
cosLookup[5694] <= 0.854640257;
cosLookup[5695] <= 0.854590471;
cosLookup[5696] <= 0.854540676;
cosLookup[5697] <= 0.854490874;
cosLookup[5698] <= 0.854441064;
cosLookup[5699] <= 0.854391246;
cosLookup[5700] <= 0.85434142;
cosLookup[5701] <= 0.854291586;
cosLookup[5702] <= 0.854241744;
cosLookup[5703] <= 0.854191895;
cosLookup[5704] <= 0.854142038;
cosLookup[5705] <= 0.854092172;
cosLookup[5706] <= 0.854042299;
cosLookup[5707] <= 0.853992419;
cosLookup[5708] <= 0.85394253;
cosLookup[5709] <= 0.853892633;
cosLookup[5710] <= 0.853842729;
cosLookup[5711] <= 0.853792817;
cosLookup[5712] <= 0.853742896;
cosLookup[5713] <= 0.853692968;
cosLookup[5714] <= 0.853643033;
cosLookup[5715] <= 0.853593089;
cosLookup[5716] <= 0.853543138;
cosLookup[5717] <= 0.853493178;
cosLookup[5718] <= 0.853443211;
cosLookup[5719] <= 0.853393236;
cosLookup[5720] <= 0.853343253;
cosLookup[5721] <= 0.853293262;
cosLookup[5722] <= 0.853243264;
cosLookup[5723] <= 0.853193257;
cosLookup[5724] <= 0.853143243;
cosLookup[5725] <= 0.853093221;
cosLookup[5726] <= 0.853043191;
cosLookup[5727] <= 0.852993153;
cosLookup[5728] <= 0.852943108;
cosLookup[5729] <= 0.852893054;
cosLookup[5730] <= 0.852842993;
cosLookup[5731] <= 0.852792924;
cosLookup[5732] <= 0.852742847;
cosLookup[5733] <= 0.852692762;
cosLookup[5734] <= 0.852642669;
cosLookup[5735] <= 0.852592569;
cosLookup[5736] <= 0.85254246;
cosLookup[5737] <= 0.852492344;
cosLookup[5738] <= 0.85244222;
cosLookup[5739] <= 0.852392088;
cosLookup[5740] <= 0.852341949;
cosLookup[5741] <= 0.852291801;
cosLookup[5742] <= 0.852241646;
cosLookup[5743] <= 0.852191483;
cosLookup[5744] <= 0.852141311;
cosLookup[5745] <= 0.852091133;
cosLookup[5746] <= 0.852040946;
cosLookup[5747] <= 0.851990751;
cosLookup[5748] <= 0.851940549;
cosLookup[5749] <= 0.851890339;
cosLookup[5750] <= 0.851840121;
cosLookup[5751] <= 0.851789895;
cosLookup[5752] <= 0.851739661;
cosLookup[5753] <= 0.85168942;
cosLookup[5754] <= 0.85163917;
cosLookup[5755] <= 0.851588913;
cosLookup[5756] <= 0.851538648;
cosLookup[5757] <= 0.851488375;
cosLookup[5758] <= 0.851438095;
cosLookup[5759] <= 0.851387806;
cosLookup[5760] <= 0.85133751;
cosLookup[5761] <= 0.851287206;
cosLookup[5762] <= 0.851236894;
cosLookup[5763] <= 0.851186574;
cosLookup[5764] <= 0.851136246;
cosLookup[5765] <= 0.851085911;
cosLookup[5766] <= 0.851035568;
cosLookup[5767] <= 0.850985217;
cosLookup[5768] <= 0.850934858;
cosLookup[5769] <= 0.850884491;
cosLookup[5770] <= 0.850834116;
cosLookup[5771] <= 0.850783734;
cosLookup[5772] <= 0.850733344;
cosLookup[5773] <= 0.850682946;
cosLookup[5774] <= 0.85063254;
cosLookup[5775] <= 0.850582126;
cosLookup[5776] <= 0.850531705;
cosLookup[5777] <= 0.850481276;
cosLookup[5778] <= 0.850430838;
cosLookup[5779] <= 0.850380393;
cosLookup[5780] <= 0.850329941;
cosLookup[5781] <= 0.85027948;
cosLookup[5782] <= 0.850229012;
cosLookup[5783] <= 0.850178536;
cosLookup[5784] <= 0.850128052;
cosLookup[5785] <= 0.85007756;
cosLookup[5786] <= 0.85002706;
cosLookup[5787] <= 0.849976553;
cosLookup[5788] <= 0.849926037;
cosLookup[5789] <= 0.849875514;
cosLookup[5790] <= 0.849824983;
cosLookup[5791] <= 0.849774445;
cosLookup[5792] <= 0.849723898;
cosLookup[5793] <= 0.849673344;
cosLookup[5794] <= 0.849622782;
cosLookup[5795] <= 0.849572212;
cosLookup[5796] <= 0.849521634;
cosLookup[5797] <= 0.849471048;
cosLookup[5798] <= 0.849420455;
cosLookup[5799] <= 0.849369854;
cosLookup[5800] <= 0.849319245;
cosLookup[5801] <= 0.849268628;
cosLookup[5802] <= 0.849218003;
cosLookup[5803] <= 0.849167371;
cosLookup[5804] <= 0.849116731;
cosLookup[5805] <= 0.849066083;
cosLookup[5806] <= 0.849015427;
cosLookup[5807] <= 0.848964763;
cosLookup[5808] <= 0.848914092;
cosLookup[5809] <= 0.848863412;
cosLookup[5810] <= 0.848812725;
cosLookup[5811] <= 0.848762031;
cosLookup[5812] <= 0.848711328;
cosLookup[5813] <= 0.848660617;
cosLookup[5814] <= 0.848609899;
cosLookup[5815] <= 0.848559173;
cosLookup[5816] <= 0.848508439;
cosLookup[5817] <= 0.848457697;
cosLookup[5818] <= 0.848406948;
cosLookup[5819] <= 0.848356191;
cosLookup[5820] <= 0.848305426;
cosLookup[5821] <= 0.848254653;
cosLookup[5822] <= 0.848203872;
cosLookup[5823] <= 0.848153084;
cosLookup[5824] <= 0.848102287;
cosLookup[5825] <= 0.848051483;
cosLookup[5826] <= 0.848000672;
cosLookup[5827] <= 0.847949852;
cosLookup[5828] <= 0.847899024;
cosLookup[5829] <= 0.847848189;
cosLookup[5830] <= 0.847797346;
cosLookup[5831] <= 0.847746495;
cosLookup[5832] <= 0.847695637;
cosLookup[5833] <= 0.84764477;
cosLookup[5834] <= 0.847593896;
cosLookup[5835] <= 0.847543014;
cosLookup[5836] <= 0.847492124;
cosLookup[5837] <= 0.847441227;
cosLookup[5838] <= 0.847390321;
cosLookup[5839] <= 0.847339408;
cosLookup[5840] <= 0.847288487;
cosLookup[5841] <= 0.847237559;
cosLookup[5842] <= 0.847186622;
cosLookup[5843] <= 0.847135678;
cosLookup[5844] <= 0.847084726;
cosLookup[5845] <= 0.847033766;
cosLookup[5846] <= 0.846982798;
cosLookup[5847] <= 0.846931823;
cosLookup[5848] <= 0.846880839;
cosLookup[5849] <= 0.846829848;
cosLookup[5850] <= 0.846778849;
cosLookup[5851] <= 0.846727843;
cosLookup[5852] <= 0.846676828;
cosLookup[5853] <= 0.846625806;
cosLookup[5854] <= 0.846574776;
cosLookup[5855] <= 0.846523739;
cosLookup[5856] <= 0.846472693;
cosLookup[5857] <= 0.84642164;
cosLookup[5858] <= 0.846370579;
cosLookup[5859] <= 0.84631951;
cosLookup[5860] <= 0.846268433;
cosLookup[5861] <= 0.846217349;
cosLookup[5862] <= 0.846166257;
cosLookup[5863] <= 0.846115157;
cosLookup[5864] <= 0.846064049;
cosLookup[5865] <= 0.846012933;
cosLookup[5866] <= 0.84596181;
cosLookup[5867] <= 0.845910679;
cosLookup[5868] <= 0.84585954;
cosLookup[5869] <= 0.845808393;
cosLookup[5870] <= 0.845757239;
cosLookup[5871] <= 0.845706077;
cosLookup[5872] <= 0.845654907;
cosLookup[5873] <= 0.845603729;
cosLookup[5874] <= 0.845552544;
cosLookup[5875] <= 0.84550135;
cosLookup[5876] <= 0.845450149;
cosLookup[5877] <= 0.84539894;
cosLookup[5878] <= 0.845347724;
cosLookup[5879] <= 0.845296499;
cosLookup[5880] <= 0.845245267;
cosLookup[5881] <= 0.845194027;
cosLookup[5882] <= 0.84514278;
cosLookup[5883] <= 0.845091524;
cosLookup[5884] <= 0.845040261;
cosLookup[5885] <= 0.84498899;
cosLookup[5886] <= 0.844937711;
cosLookup[5887] <= 0.844886425;
cosLookup[5888] <= 0.84483513;
cosLookup[5889] <= 0.844783828;
cosLookup[5890] <= 0.844732519;
cosLookup[5891] <= 0.844681201;
cosLookup[5892] <= 0.844629876;
cosLookup[5893] <= 0.844578543;
cosLookup[5894] <= 0.844527202;
cosLookup[5895] <= 0.844475853;
cosLookup[5896] <= 0.844424497;
cosLookup[5897] <= 0.844373132;
cosLookup[5898] <= 0.84432176;
cosLookup[5899] <= 0.844270381;
cosLookup[5900] <= 0.844218993;
cosLookup[5901] <= 0.844167598;
cosLookup[5902] <= 0.844116195;
cosLookup[5903] <= 0.844064784;
cosLookup[5904] <= 0.844013366;
cosLookup[5905] <= 0.84396194;
cosLookup[5906] <= 0.843910506;
cosLookup[5907] <= 0.843859064;
cosLookup[5908] <= 0.843807614;
cosLookup[5909] <= 0.843756157;
cosLookup[5910] <= 0.843704692;
cosLookup[5911] <= 0.843653219;
cosLookup[5912] <= 0.843601739;
cosLookup[5913] <= 0.84355025;
cosLookup[5914] <= 0.843498754;
cosLookup[5915] <= 0.84344725;
cosLookup[5916] <= 0.843395739;
cosLookup[5917] <= 0.843344219;
cosLookup[5918] <= 0.843292692;
cosLookup[5919] <= 0.843241158;
cosLookup[5920] <= 0.843189615;
cosLookup[5921] <= 0.843138065;
cosLookup[5922] <= 0.843086507;
cosLookup[5923] <= 0.843034941;
cosLookup[5924] <= 0.842983367;
cosLookup[5925] <= 0.842931786;
cosLookup[5926] <= 0.842880197;
cosLookup[5927] <= 0.8428286;
cosLookup[5928] <= 0.842776995;
cosLookup[5929] <= 0.842725383;
cosLookup[5930] <= 0.842673763;
cosLookup[5931] <= 0.842622135;
cosLookup[5932] <= 0.842570499;
cosLookup[5933] <= 0.842518856;
cosLookup[5934] <= 0.842467205;
cosLookup[5935] <= 0.842415546;
cosLookup[5936] <= 0.84236388;
cosLookup[5937] <= 0.842312205;
cosLookup[5938] <= 0.842260523;
cosLookup[5939] <= 0.842208834;
cosLookup[5940] <= 0.842157136;
cosLookup[5941] <= 0.842105431;
cosLookup[5942] <= 0.842053718;
cosLookup[5943] <= 0.842001997;
cosLookup[5944] <= 0.841950269;
cosLookup[5945] <= 0.841898532;
cosLookup[5946] <= 0.841846788;
cosLookup[5947] <= 0.841795037;
cosLookup[5948] <= 0.841743277;
cosLookup[5949] <= 0.84169151;
cosLookup[5950] <= 0.841639735;
cosLookup[5951] <= 0.841587952;
cosLookup[5952] <= 0.841536162;
cosLookup[5953] <= 0.841484364;
cosLookup[5954] <= 0.841432558;
cosLookup[5955] <= 0.841380744;
cosLookup[5956] <= 0.841328923;
cosLookup[5957] <= 0.841277094;
cosLookup[5958] <= 0.841225257;
cosLookup[5959] <= 0.841173413;
cosLookup[5960] <= 0.84112156;
cosLookup[5961] <= 0.8410697;
cosLookup[5962] <= 0.841017833;
cosLookup[5963] <= 0.840965957;
cosLookup[5964] <= 0.840914074;
cosLookup[5965] <= 0.840862183;
cosLookup[5966] <= 0.840810284;
cosLookup[5967] <= 0.840758378;
cosLookup[5968] <= 0.840706464;
cosLookup[5969] <= 0.840654542;
cosLookup[5970] <= 0.840602613;
cosLookup[5971] <= 0.840550675;
cosLookup[5972] <= 0.84049873;
cosLookup[5973] <= 0.840446777;
cosLookup[5974] <= 0.840394817;
cosLookup[5975] <= 0.840342849;
cosLookup[5976] <= 0.840290873;
cosLookup[5977] <= 0.840238889;
cosLookup[5978] <= 0.840186898;
cosLookup[5979] <= 0.840134899;
cosLookup[5980] <= 0.840082892;
cosLookup[5981] <= 0.840030877;
cosLookup[5982] <= 0.839978855;
cosLookup[5983] <= 0.839926825;
cosLookup[5984] <= 0.839874787;
cosLookup[5985] <= 0.839822742;
cosLookup[5986] <= 0.839770689;
cosLookup[5987] <= 0.839718628;
cosLookup[5988] <= 0.839666559;
cosLookup[5989] <= 0.839614483;
cosLookup[5990] <= 0.839562399;
cosLookup[5991] <= 0.839510307;
cosLookup[5992] <= 0.839458208;
cosLookup[5993] <= 0.839406101;
cosLookup[5994] <= 0.839353986;
cosLookup[5995] <= 0.839301863;
cosLookup[5996] <= 0.839249733;
cosLookup[5997] <= 0.839197595;
cosLookup[5998] <= 0.839145449;
cosLookup[5999] <= 0.839093295;
cosLookup[6000] <= 0.839041134;
cosLookup[6001] <= 0.838988965;
cosLookup[6002] <= 0.838936789;
cosLookup[6003] <= 0.838884604;
cosLookup[6004] <= 0.838832412;
cosLookup[6005] <= 0.838780213;
cosLookup[6006] <= 0.838728005;
cosLookup[6007] <= 0.83867579;
cosLookup[6008] <= 0.838623567;
cosLookup[6009] <= 0.838571336;
cosLookup[6010] <= 0.838519098;
cosLookup[6011] <= 0.838466852;
cosLookup[6012] <= 0.838414598;
cosLookup[6013] <= 0.838362337;
cosLookup[6014] <= 0.838310068;
cosLookup[6015] <= 0.838257791;
cosLookup[6016] <= 0.838205506;
cosLookup[6017] <= 0.838153214;
cosLookup[6018] <= 0.838100914;
cosLookup[6019] <= 0.838048607;
cosLookup[6020] <= 0.837996291;
cosLookup[6021] <= 0.837943968;
cosLookup[6022] <= 0.837891637;
cosLookup[6023] <= 0.837839299;
cosLookup[6024] <= 0.837786953;
cosLookup[6025] <= 0.837734599;
cosLookup[6026] <= 0.837682237;
cosLookup[6027] <= 0.837629868;
cosLookup[6028] <= 0.837577491;
cosLookup[6029] <= 0.837525106;
cosLookup[6030] <= 0.837472714;
cosLookup[6031] <= 0.837420314;
cosLookup[6032] <= 0.837367906;
cosLookup[6033] <= 0.837315491;
cosLookup[6034] <= 0.837263067;
cosLookup[6035] <= 0.837210637;
cosLookup[6036] <= 0.837158198;
cosLookup[6037] <= 0.837105752;
cosLookup[6038] <= 0.837053298;
cosLookup[6039] <= 0.837000836;
cosLookup[6040] <= 0.836948367;
cosLookup[6041] <= 0.83689589;
cosLookup[6042] <= 0.836843405;
cosLookup[6043] <= 0.836790913;
cosLookup[6044] <= 0.836738412;
cosLookup[6045] <= 0.836685905;
cosLookup[6046] <= 0.836633389;
cosLookup[6047] <= 0.836580866;
cosLookup[6048] <= 0.836528335;
cosLookup[6049] <= 0.836475796;
cosLookup[6050] <= 0.83642325;
cosLookup[6051] <= 0.836370696;
cosLookup[6052] <= 0.836318135;
cosLookup[6053] <= 0.836265565;
cosLookup[6054] <= 0.836212988;
cosLookup[6055] <= 0.836160404;
cosLookup[6056] <= 0.836107811;
cosLookup[6057] <= 0.836055211;
cosLookup[6058] <= 0.836002603;
cosLookup[6059] <= 0.835949988;
cosLookup[6060] <= 0.835897365;
cosLookup[6061] <= 0.835844734;
cosLookup[6062] <= 0.835792095;
cosLookup[6063] <= 0.835739449;
cosLookup[6064] <= 0.835686795;
cosLookup[6065] <= 0.835634134;
cosLookup[6066] <= 0.835581465;
cosLookup[6067] <= 0.835528788;
cosLookup[6068] <= 0.835476103;
cosLookup[6069] <= 0.835423411;
cosLookup[6070] <= 0.835370711;
cosLookup[6071] <= 0.835318003;
cosLookup[6072] <= 0.835265288;
cosLookup[6073] <= 0.835212565;
cosLookup[6074] <= 0.835159834;
cosLookup[6075] <= 0.835107096;
cosLookup[6076] <= 0.83505435;
cosLookup[6077] <= 0.835001596;
cosLookup[6078] <= 0.834948835;
cosLookup[6079] <= 0.834896066;
cosLookup[6080] <= 0.834843289;
cosLookup[6081] <= 0.834790505;
cosLookup[6082] <= 0.834737712;
cosLookup[6083] <= 0.834684913;
cosLookup[6084] <= 0.834632105;
cosLookup[6085] <= 0.83457929;
cosLookup[6086] <= 0.834526467;
cosLookup[6087] <= 0.834473637;
cosLookup[6088] <= 0.834420799;
cosLookup[6089] <= 0.834367953;
cosLookup[6090] <= 0.8343151;
cosLookup[6091] <= 0.834262239;
cosLookup[6092] <= 0.83420937;
cosLookup[6093] <= 0.834156493;
cosLookup[6094] <= 0.834103609;
cosLookup[6095] <= 0.834050717;
cosLookup[6096] <= 0.833997818;
cosLookup[6097] <= 0.833944911;
cosLookup[6098] <= 0.833891996;
cosLookup[6099] <= 0.833839073;
cosLookup[6100] <= 0.833786143;
cosLookup[6101] <= 0.833733206;
cosLookup[6102] <= 0.83368026;
cosLookup[6103] <= 0.833627307;
cosLookup[6104] <= 0.833574346;
cosLookup[6105] <= 0.833521378;
cosLookup[6106] <= 0.833468402;
cosLookup[6107] <= 0.833415418;
cosLookup[6108] <= 0.833362426;
cosLookup[6109] <= 0.833309427;
cosLookup[6110] <= 0.833256421;
cosLookup[6111] <= 0.833203406;
cosLookup[6112] <= 0.833150384;
cosLookup[6113] <= 0.833097354;
cosLookup[6114] <= 0.833044317;
cosLookup[6115] <= 0.832991272;
cosLookup[6116] <= 0.832938219;
cosLookup[6117] <= 0.832885159;
cosLookup[6118] <= 0.832832091;
cosLookup[6119] <= 0.832779015;
cosLookup[6120] <= 0.832725932;
cosLookup[6121] <= 0.832672841;
cosLookup[6122] <= 0.832619742;
cosLookup[6123] <= 0.832566636;
cosLookup[6124] <= 0.832513522;
cosLookup[6125] <= 0.8324604;
cosLookup[6126] <= 0.832407271;
cosLookup[6127] <= 0.832354134;
cosLookup[6128] <= 0.83230099;
cosLookup[6129] <= 0.832247837;
cosLookup[6130] <= 0.832194677;
cosLookup[6131] <= 0.83214151;
cosLookup[6132] <= 0.832088335;
cosLookup[6133] <= 0.832035152;
cosLookup[6134] <= 0.831981962;
cosLookup[6135] <= 0.831928763;
cosLookup[6136] <= 0.831875558;
cosLookup[6137] <= 0.831822344;
cosLookup[6138] <= 0.831769123;
cosLookup[6139] <= 0.831715894;
cosLookup[6140] <= 0.831662658;
cosLookup[6141] <= 0.831609414;
cosLookup[6142] <= 0.831556163;
cosLookup[6143] <= 0.831502903;
cosLookup[6144] <= 0.831449636;
cosLookup[6145] <= 0.831396362;
cosLookup[6146] <= 0.83134308;
cosLookup[6147] <= 0.83128979;
cosLookup[6148] <= 0.831236492;
cosLookup[6149] <= 0.831183187;
cosLookup[6150] <= 0.831129874;
cosLookup[6151] <= 0.831076554;
cosLookup[6152] <= 0.831023226;
cosLookup[6153] <= 0.83096989;
cosLookup[6154] <= 0.830916547;
cosLookup[6155] <= 0.830863196;
cosLookup[6156] <= 0.830809837;
cosLookup[6157] <= 0.830756471;
cosLookup[6158] <= 0.830703097;
cosLookup[6159] <= 0.830649716;
cosLookup[6160] <= 0.830596326;
cosLookup[6161] <= 0.83054293;
cosLookup[6162] <= 0.830489525;
cosLookup[6163] <= 0.830436113;
cosLookup[6164] <= 0.830382693;
cosLookup[6165] <= 0.830329266;
cosLookup[6166] <= 0.830275831;
cosLookup[6167] <= 0.830222388;
cosLookup[6168] <= 0.830168938;
cosLookup[6169] <= 0.83011548;
cosLookup[6170] <= 0.830062015;
cosLookup[6171] <= 0.830008542;
cosLookup[6172] <= 0.829955061;
cosLookup[6173] <= 0.829901573;
cosLookup[6174] <= 0.829848077;
cosLookup[6175] <= 0.829794573;
cosLookup[6176] <= 0.829741062;
cosLookup[6177] <= 0.829687543;
cosLookup[6178] <= 0.829634016;
cosLookup[6179] <= 0.829580482;
cosLookup[6180] <= 0.82952694;
cosLookup[6181] <= 0.829473391;
cosLookup[6182] <= 0.829419834;
cosLookup[6183] <= 0.829366269;
cosLookup[6184] <= 0.829312697;
cosLookup[6185] <= 0.829259117;
cosLookup[6186] <= 0.829205529;
cosLookup[6187] <= 0.829151934;
cosLookup[6188] <= 0.829098332;
cosLookup[6189] <= 0.829044721;
cosLookup[6190] <= 0.828991103;
cosLookup[6191] <= 0.828937478;
cosLookup[6192] <= 0.828883844;
cosLookup[6193] <= 0.828830203;
cosLookup[6194] <= 0.828776555;
cosLookup[6195] <= 0.828722899;
cosLookup[6196] <= 0.828669235;
cosLookup[6197] <= 0.828615564;
cosLookup[6198] <= 0.828561885;
cosLookup[6199] <= 0.828508198;
cosLookup[6200] <= 0.828454504;
cosLookup[6201] <= 0.828400802;
cosLookup[6202] <= 0.828347093;
cosLookup[6203] <= 0.828293376;
cosLookup[6204] <= 0.828239651;
cosLookup[6205] <= 0.828185919;
cosLookup[6206] <= 0.828132179;
cosLookup[6207] <= 0.828078431;
cosLookup[6208] <= 0.828024676;
cosLookup[6209] <= 0.827970913;
cosLookup[6210] <= 0.827917143;
cosLookup[6211] <= 0.827863365;
cosLookup[6212] <= 0.82780958;
cosLookup[6213] <= 0.827755786;
cosLookup[6214] <= 0.827701986;
cosLookup[6215] <= 0.827648177;
cosLookup[6216] <= 0.827594361;
cosLookup[6217] <= 0.827540538;
cosLookup[6218] <= 0.827486706;
cosLookup[6219] <= 0.827432868;
cosLookup[6220] <= 0.827379021;
cosLookup[6221] <= 0.827325167;
cosLookup[6222] <= 0.827271306;
cosLookup[6223] <= 0.827217436;
cosLookup[6224] <= 0.827163559;
cosLookup[6225] <= 0.827109675;
cosLookup[6226] <= 0.827055783;
cosLookup[6227] <= 0.827001883;
cosLookup[6228] <= 0.826947976;
cosLookup[6229] <= 0.826894061;
cosLookup[6230] <= 0.826840139;
cosLookup[6231] <= 0.826786209;
cosLookup[6232] <= 0.826732271;
cosLookup[6233] <= 0.826678326;
cosLookup[6234] <= 0.826624373;
cosLookup[6235] <= 0.826570412;
cosLookup[6236] <= 0.826516444;
cosLookup[6237] <= 0.826462469;
cosLookup[6238] <= 0.826408485;
cosLookup[6239] <= 0.826354495;
cosLookup[6240] <= 0.826300496;
cosLookup[6241] <= 0.82624649;
cosLookup[6242] <= 0.826192476;
cosLookup[6243] <= 0.826138455;
cosLookup[6244] <= 0.826084426;
cosLookup[6245] <= 0.82603039;
cosLookup[6246] <= 0.825976346;
cosLookup[6247] <= 0.825922294;
cosLookup[6248] <= 0.825868235;
cosLookup[6249] <= 0.825814168;
cosLookup[6250] <= 0.825760094;
cosLookup[6251] <= 0.825706012;
cosLookup[6252] <= 0.825651922;
cosLookup[6253] <= 0.825597825;
cosLookup[6254] <= 0.82554372;
cosLookup[6255] <= 0.825489608;
cosLookup[6256] <= 0.825435488;
cosLookup[6257] <= 0.825381361;
cosLookup[6258] <= 0.825327226;
cosLookup[6259] <= 0.825273083;
cosLookup[6260] <= 0.825218933;
cosLookup[6261] <= 0.825164775;
cosLookup[6262] <= 0.825110609;
cosLookup[6263] <= 0.825056436;
cosLookup[6264] <= 0.825002256;
cosLookup[6265] <= 0.824948067;
cosLookup[6266] <= 0.824893872;
cosLookup[6267] <= 0.824839668;
cosLookup[6268] <= 0.824785457;
cosLookup[6269] <= 0.824731239;
cosLookup[6270] <= 0.824677013;
cosLookup[6271] <= 0.824622779;
cosLookup[6272] <= 0.824568538;
cosLookup[6273] <= 0.824514289;
cosLookup[6274] <= 0.824460032;
cosLookup[6275] <= 0.824405768;
cosLookup[6276] <= 0.824351497;
cosLookup[6277] <= 0.824297218;
cosLookup[6278] <= 0.824242931;
cosLookup[6279] <= 0.824188636;
cosLookup[6280] <= 0.824134335;
cosLookup[6281] <= 0.824080025;
cosLookup[6282] <= 0.824025708;
cosLookup[6283] <= 0.823971383;
cosLookup[6284] <= 0.823917051;
cosLookup[6285] <= 0.823862711;
cosLookup[6286] <= 0.823808364;
cosLookup[6287] <= 0.823754009;
cosLookup[6288] <= 0.823699647;
cosLookup[6289] <= 0.823645277;
cosLookup[6290] <= 0.823590899;
cosLookup[6291] <= 0.823536514;
cosLookup[6292] <= 0.823482121;
cosLookup[6293] <= 0.823427721;
cosLookup[6294] <= 0.823373313;
cosLookup[6295] <= 0.823318897;
cosLookup[6296] <= 0.823264474;
cosLookup[6297] <= 0.823210043;
cosLookup[6298] <= 0.823155605;
cosLookup[6299] <= 0.823101159;
cosLookup[6300] <= 0.823046706;
cosLookup[6301] <= 0.822992245;
cosLookup[6302] <= 0.822937777;
cosLookup[6303] <= 0.822883301;
cosLookup[6304] <= 0.822828817;
cosLookup[6305] <= 0.822774326;
cosLookup[6306] <= 0.822719827;
cosLookup[6307] <= 0.822665321;
cosLookup[6308] <= 0.822610807;
cosLookup[6309] <= 0.822556286;
cosLookup[6310] <= 0.822501757;
cosLookup[6311] <= 0.82244722;
cosLookup[6312] <= 0.822392676;
cosLookup[6313] <= 0.822338124;
cosLookup[6314] <= 0.822283565;
cosLookup[6315] <= 0.822228998;
cosLookup[6316] <= 0.822174424;
cosLookup[6317] <= 0.822119842;
cosLookup[6318] <= 0.822065253;
cosLookup[6319] <= 0.822010656;
cosLookup[6320] <= 0.821956051;
cosLookup[6321] <= 0.821901439;
cosLookup[6322] <= 0.821846819;
cosLookup[6323] <= 0.821792192;
cosLookup[6324] <= 0.821737557;
cosLookup[6325] <= 0.821682915;
cosLookup[6326] <= 0.821628265;
cosLookup[6327] <= 0.821573608;
cosLookup[6328] <= 0.821518943;
cosLookup[6329] <= 0.82146427;
cosLookup[6330] <= 0.82140959;
cosLookup[6331] <= 0.821354902;
cosLookup[6332] <= 0.821300207;
cosLookup[6333] <= 0.821245504;
cosLookup[6334] <= 0.821190794;
cosLookup[6335] <= 0.821136076;
cosLookup[6336] <= 0.821081351;
cosLookup[6337] <= 0.821026618;
cosLookup[6338] <= 0.820971877;
cosLookup[6339] <= 0.820917129;
cosLookup[6340] <= 0.820862374;
cosLookup[6341] <= 0.820807611;
cosLookup[6342] <= 0.82075284;
cosLookup[6343] <= 0.820698062;
cosLookup[6344] <= 0.820643276;
cosLookup[6345] <= 0.820588483;
cosLookup[6346] <= 0.820533682;
cosLookup[6347] <= 0.820478873;
cosLookup[6348] <= 0.820424057;
cosLookup[6349] <= 0.820369234;
cosLookup[6350] <= 0.820314403;
cosLookup[6351] <= 0.820259564;
cosLookup[6352] <= 0.820204718;
cosLookup[6353] <= 0.820149864;
cosLookup[6354] <= 0.820095003;
cosLookup[6355] <= 0.820040135;
cosLookup[6356] <= 0.819985258;
cosLookup[6357] <= 0.819930374;
cosLookup[6358] <= 0.819875483;
cosLookup[6359] <= 0.819820584;
cosLookup[6360] <= 0.819765678;
cosLookup[6361] <= 0.819710764;
cosLookup[6362] <= 0.819655842;
cosLookup[6363] <= 0.819600913;
cosLookup[6364] <= 0.819545977;
cosLookup[6365] <= 0.819491033;
cosLookup[6366] <= 0.819436081;
cosLookup[6367] <= 0.819381122;
cosLookup[6368] <= 0.819326155;
cosLookup[6369] <= 0.819271181;
cosLookup[6370] <= 0.819216199;
cosLookup[6371] <= 0.81916121;
cosLookup[6372] <= 0.819106213;
cosLookup[6373] <= 0.819051209;
cosLookup[6374] <= 0.818996197;
cosLookup[6375] <= 0.818941177;
cosLookup[6376] <= 0.818886151;
cosLookup[6377] <= 0.818831116;
cosLookup[6378] <= 0.818776074;
cosLookup[6379] <= 0.818721025;
cosLookup[6380] <= 0.818665967;
cosLookup[6381] <= 0.818610903;
cosLookup[6382] <= 0.818555831;
cosLookup[6383] <= 0.818500751;
cosLookup[6384] <= 0.818445664;
cosLookup[6385] <= 0.818390569;
cosLookup[6386] <= 0.818335467;
cosLookup[6387] <= 0.818280357;
cosLookup[6388] <= 0.81822524;
cosLookup[6389] <= 0.818170115;
cosLookup[6390] <= 0.818114983;
cosLookup[6391] <= 0.818059843;
cosLookup[6392] <= 0.818004696;
cosLookup[6393] <= 0.817949541;
cosLookup[6394] <= 0.817894379;
cosLookup[6395] <= 0.817839209;
cosLookup[6396] <= 0.817784032;
cosLookup[6397] <= 0.817728847;
cosLookup[6398] <= 0.817673654;
cosLookup[6399] <= 0.817618454;
cosLookup[6400] <= 0.817563247;
cosLookup[6401] <= 0.817508032;
cosLookup[6402] <= 0.817452809;
cosLookup[6403] <= 0.817397579;
cosLookup[6404] <= 0.817342342;
cosLookup[6405] <= 0.817287097;
cosLookup[6406] <= 0.817231844;
cosLookup[6407] <= 0.817176584;
cosLookup[6408] <= 0.817121317;
cosLookup[6409] <= 0.817066041;
cosLookup[6410] <= 0.817010759;
cosLookup[6411] <= 0.816955469;
cosLookup[6412] <= 0.816900171;
cosLookup[6413] <= 0.816844866;
cosLookup[6414] <= 0.816789553;
cosLookup[6415] <= 0.816734233;
cosLookup[6416] <= 0.816678906;
cosLookup[6417] <= 0.81662357;
cosLookup[6418] <= 0.816568228;
cosLookup[6419] <= 0.816512878;
cosLookup[6420] <= 0.81645752;
cosLookup[6421] <= 0.816402155;
cosLookup[6422] <= 0.816346782;
cosLookup[6423] <= 0.816291402;
cosLookup[6424] <= 0.816236014;
cosLookup[6425] <= 0.816180619;
cosLookup[6426] <= 0.816125216;
cosLookup[6427] <= 0.816069806;
cosLookup[6428] <= 0.816014388;
cosLookup[6429] <= 0.815958963;
cosLookup[6430] <= 0.81590353;
cosLookup[6431] <= 0.81584809;
cosLookup[6432] <= 0.815792642;
cosLookup[6433] <= 0.815737187;
cosLookup[6434] <= 0.815681724;
cosLookup[6435] <= 0.815626254;
cosLookup[6436] <= 0.815570776;
cosLookup[6437] <= 0.815515291;
cosLookup[6438] <= 0.815459799;
cosLookup[6439] <= 0.815404298;
cosLookup[6440] <= 0.815348791;
cosLookup[6441] <= 0.815293275;
cosLookup[6442] <= 0.815237753;
cosLookup[6443] <= 0.815182223;
cosLookup[6444] <= 0.815126685;
cosLookup[6445] <= 0.81507114;
cosLookup[6446] <= 0.815015587;
cosLookup[6447] <= 0.814960027;
cosLookup[6448] <= 0.814904459;
cosLookup[6449] <= 0.814848884;
cosLookup[6450] <= 0.814793301;
cosLookup[6451] <= 0.814737711;
cosLookup[6452] <= 0.814682114;
cosLookup[6453] <= 0.814626509;
cosLookup[6454] <= 0.814570896;
cosLookup[6455] <= 0.814515276;
cosLookup[6456] <= 0.814459648;
cosLookup[6457] <= 0.814404013;
cosLookup[6458] <= 0.814348371;
cosLookup[6459] <= 0.814292721;
cosLookup[6460] <= 0.814237063;
cosLookup[6461] <= 0.814181398;
cosLookup[6462] <= 0.814125726;
cosLookup[6463] <= 0.814070046;
cosLookup[6464] <= 0.814014358;
cosLookup[6465] <= 0.813958663;
cosLookup[6466] <= 0.813902961;
cosLookup[6467] <= 0.813847251;
cosLookup[6468] <= 0.813791534;
cosLookup[6469] <= 0.813735809;
cosLookup[6470] <= 0.813680077;
cosLookup[6471] <= 0.813624337;
cosLookup[6472] <= 0.813568589;
cosLookup[6473] <= 0.813512835;
cosLookup[6474] <= 0.813457072;
cosLookup[6475] <= 0.813401303;
cosLookup[6476] <= 0.813345525;
cosLookup[6477] <= 0.813289741;
cosLookup[6478] <= 0.813233949;
cosLookup[6479] <= 0.813178149;
cosLookup[6480] <= 0.813122342;
cosLookup[6481] <= 0.813066527;
cosLookup[6482] <= 0.813010705;
cosLookup[6483] <= 0.812954876;
cosLookup[6484] <= 0.812899039;
cosLookup[6485] <= 0.812843194;
cosLookup[6486] <= 0.812787342;
cosLookup[6487] <= 0.812731483;
cosLookup[6488] <= 0.812675616;
cosLookup[6489] <= 0.812619741;
cosLookup[6490] <= 0.81256386;
cosLookup[6491] <= 0.81250797;
cosLookup[6492] <= 0.812452073;
cosLookup[6493] <= 0.812396169;
cosLookup[6494] <= 0.812340257;
cosLookup[6495] <= 0.812284338;
cosLookup[6496] <= 0.812228412;
cosLookup[6497] <= 0.812172478;
cosLookup[6498] <= 0.812116536;
cosLookup[6499] <= 0.812060587;
cosLookup[6500] <= 0.81200463;
cosLookup[6501] <= 0.811948666;
cosLookup[6502] <= 0.811892695;
cosLookup[6503] <= 0.811836716;
cosLookup[6504] <= 0.81178073;
cosLookup[6505] <= 0.811724736;
cosLookup[6506] <= 0.811668734;
cosLookup[6507] <= 0.811612726;
cosLookup[6508] <= 0.81155671;
cosLookup[6509] <= 0.811500686;
cosLookup[6510] <= 0.811444655;
cosLookup[6511] <= 0.811388616;
cosLookup[6512] <= 0.81133257;
cosLookup[6513] <= 0.811276516;
cosLookup[6514] <= 0.811220456;
cosLookup[6515] <= 0.811164387;
cosLookup[6516] <= 0.811108311;
cosLookup[6517] <= 0.811052228;
cosLookup[6518] <= 0.810996137;
cosLookup[6519] <= 0.810940039;
cosLookup[6520] <= 0.810883933;
cosLookup[6521] <= 0.81082782;
cosLookup[6522] <= 0.810771699;
cosLookup[6523] <= 0.810715571;
cosLookup[6524] <= 0.810659436;
cosLookup[6525] <= 0.810603293;
cosLookup[6526] <= 0.810547142;
cosLookup[6527] <= 0.810490984;
cosLookup[6528] <= 0.810434819;
cosLookup[6529] <= 0.810378646;
cosLookup[6530] <= 0.810322466;
cosLookup[6531] <= 0.810266278;
cosLookup[6532] <= 0.810210083;
cosLookup[6533] <= 0.810153881;
cosLookup[6534] <= 0.810097671;
cosLookup[6535] <= 0.810041453;
cosLookup[6536] <= 0.809985228;
cosLookup[6537] <= 0.809928996;
cosLookup[6538] <= 0.809872756;
cosLookup[6539] <= 0.809816509;
cosLookup[6540] <= 0.809760254;
cosLookup[6541] <= 0.809703992;
cosLookup[6542] <= 0.809647722;
cosLookup[6543] <= 0.809591445;
cosLookup[6544] <= 0.809535161;
cosLookup[6545] <= 0.809478869;
cosLookup[6546] <= 0.809422569;
cosLookup[6547] <= 0.809366263;
cosLookup[6548] <= 0.809309948;
cosLookup[6549] <= 0.809253627;
cosLookup[6550] <= 0.809197298;
cosLookup[6551] <= 0.809140961;
cosLookup[6552] <= 0.809084617;
cosLookup[6553] <= 0.809028266;
cosLookup[6554] <= 0.808971907;
cosLookup[6555] <= 0.80891554;
cosLookup[6556] <= 0.808859167;
cosLookup[6557] <= 0.808802785;
cosLookup[6558] <= 0.808746397;
cosLookup[6559] <= 0.808690001;
cosLookup[6560] <= 0.808633597;
cosLookup[6561] <= 0.808577186;
cosLookup[6562] <= 0.808520768;
cosLookup[6563] <= 0.808464342;
cosLookup[6564] <= 0.808407909;
cosLookup[6565] <= 0.808351468;
cosLookup[6566] <= 0.80829502;
cosLookup[6567] <= 0.808238565;
cosLookup[6568] <= 0.808182102;
cosLookup[6569] <= 0.808125631;
cosLookup[6570] <= 0.808069154;
cosLookup[6571] <= 0.808012668;
cosLookup[6572] <= 0.807956176;
cosLookup[6573] <= 0.807899676;
cosLookup[6574] <= 0.807843168;
cosLookup[6575] <= 0.807786653;
cosLookup[6576] <= 0.807730131;
cosLookup[6577] <= 0.807673601;
cosLookup[6578] <= 0.807617064;
cosLookup[6579] <= 0.807560519;
cosLookup[6580] <= 0.807503967;
cosLookup[6581] <= 0.807447408;
cosLookup[6582] <= 0.807390841;
cosLookup[6583] <= 0.807334266;
cosLookup[6584] <= 0.807277685;
cosLookup[6585] <= 0.807221095;
cosLookup[6586] <= 0.807164499;
cosLookup[6587] <= 0.807107895;
cosLookup[6588] <= 0.807051283;
cosLookup[6589] <= 0.806994665;
cosLookup[6590] <= 0.806938038;
cosLookup[6591] <= 0.806881405;
cosLookup[6592] <= 0.806824763;
cosLookup[6593] <= 0.806768115;
cosLookup[6594] <= 0.806711459;
cosLookup[6595] <= 0.806654796;
cosLookup[6596] <= 0.806598125;
cosLookup[6597] <= 0.806541447;
cosLookup[6598] <= 0.806484761;
cosLookup[6599] <= 0.806428068;
cosLookup[6600] <= 0.806371368;
cosLookup[6601] <= 0.80631466;
cosLookup[6602] <= 0.806257945;
cosLookup[6603] <= 0.806201222;
cosLookup[6604] <= 0.806144492;
cosLookup[6605] <= 0.806087754;
cosLookup[6606] <= 0.806031009;
cosLookup[6607] <= 0.805974257;
cosLookup[6608] <= 0.805917497;
cosLookup[6609] <= 0.80586073;
cosLookup[6610] <= 0.805803956;
cosLookup[6611] <= 0.805747174;
cosLookup[6612] <= 0.805690384;
cosLookup[6613] <= 0.805633588;
cosLookup[6614] <= 0.805576783;
cosLookup[6615] <= 0.805519972;
cosLookup[6616] <= 0.805463153;
cosLookup[6617] <= 0.805406327;
cosLookup[6618] <= 0.805349493;
cosLookup[6619] <= 0.805292652;
cosLookup[6620] <= 0.805235803;
cosLookup[6621] <= 0.805178947;
cosLookup[6622] <= 0.805122084;
cosLookup[6623] <= 0.805065213;
cosLookup[6624] <= 0.805008335;
cosLookup[6625] <= 0.804951449;
cosLookup[6626] <= 0.804894556;
cosLookup[6627] <= 0.804837656;
cosLookup[6628] <= 0.804780748;
cosLookup[6629] <= 0.804723833;
cosLookup[6630] <= 0.80466691;
cosLookup[6631] <= 0.80460998;
cosLookup[6632] <= 0.804553043;
cosLookup[6633] <= 0.804496098;
cosLookup[6634] <= 0.804439146;
cosLookup[6635] <= 0.804382186;
cosLookup[6636] <= 0.804325219;
cosLookup[6637] <= 0.804268245;
cosLookup[6638] <= 0.804211263;
cosLookup[6639] <= 0.804154274;
cosLookup[6640] <= 0.804097277;
cosLookup[6641] <= 0.804040273;
cosLookup[6642] <= 0.803983262;
cosLookup[6643] <= 0.803926243;
cosLookup[6644] <= 0.803869217;
cosLookup[6645] <= 0.803812184;
cosLookup[6646] <= 0.803755143;
cosLookup[6647] <= 0.803698095;
cosLookup[6648] <= 0.803641039;
cosLookup[6649] <= 0.803583976;
cosLookup[6650] <= 0.803526905;
cosLookup[6651] <= 0.803469828;
cosLookup[6652] <= 0.803412742;
cosLookup[6653] <= 0.80335565;
cosLookup[6654] <= 0.80329855;
cosLookup[6655] <= 0.803241442;
cosLookup[6656] <= 0.803184328;
cosLookup[6657] <= 0.803127206;
cosLookup[6658] <= 0.803070076;
cosLookup[6659] <= 0.803012939;
cosLookup[6660] <= 0.802955795;
cosLookup[6661] <= 0.802898643;
cosLookup[6662] <= 0.802841484;
cosLookup[6663] <= 0.802784318;
cosLookup[6664] <= 0.802727144;
cosLookup[6665] <= 0.802669963;
cosLookup[6666] <= 0.802612774;
cosLookup[6667] <= 0.802555578;
cosLookup[6668] <= 0.802498375;
cosLookup[6669] <= 0.802441164;
cosLookup[6670] <= 0.802383946;
cosLookup[6671] <= 0.802326721;
cosLookup[6672] <= 0.802269488;
cosLookup[6673] <= 0.802212248;
cosLookup[6674] <= 0.802155;
cosLookup[6675] <= 0.802097745;
cosLookup[6676] <= 0.802040483;
cosLookup[6677] <= 0.801983213;
cosLookup[6678] <= 0.801925936;
cosLookup[6679] <= 0.801868652;
cosLookup[6680] <= 0.80181136;
cosLookup[6681] <= 0.801754061;
cosLookup[6682] <= 0.801696754;
cosLookup[6683] <= 0.80163944;
cosLookup[6684] <= 0.801582119;
cosLookup[6685] <= 0.80152479;
cosLookup[6686] <= 0.801467454;
cosLookup[6687] <= 0.801410111;
cosLookup[6688] <= 0.80135276;
cosLookup[6689] <= 0.801295402;
cosLookup[6690] <= 0.801238036;
cosLookup[6691] <= 0.801180664;
cosLookup[6692] <= 0.801123283;
cosLookup[6693] <= 0.801065896;
cosLookup[6694] <= 0.801008501;
cosLookup[6695] <= 0.800951098;
cosLookup[6696] <= 0.800893689;
cosLookup[6697] <= 0.800836272;
cosLookup[6698] <= 0.800778847;
cosLookup[6699] <= 0.800721416;
cosLookup[6700] <= 0.800663976;
cosLookup[6701] <= 0.80060653;
cosLookup[6702] <= 0.800549076;
cosLookup[6703] <= 0.800491615;
cosLookup[6704] <= 0.800434146;
cosLookup[6705] <= 0.80037667;
cosLookup[6706] <= 0.800319187;
cosLookup[6707] <= 0.800261696;
cosLookup[6708] <= 0.800204198;
cosLookup[6709] <= 0.800146693;
cosLookup[6710] <= 0.80008918;
cosLookup[6711] <= 0.80003166;
cosLookup[6712] <= 0.799974133;
cosLookup[6713] <= 0.799916598;
cosLookup[6714] <= 0.799859056;
cosLookup[6715] <= 0.799801507;
cosLookup[6716] <= 0.79974395;
cosLookup[6717] <= 0.799686386;
cosLookup[6718] <= 0.799628814;
cosLookup[6719] <= 0.799571235;
cosLookup[6720] <= 0.799513649;
cosLookup[6721] <= 0.799456055;
cosLookup[6722] <= 0.799398454;
cosLookup[6723] <= 0.799340846;
cosLookup[6724] <= 0.79928323;
cosLookup[6725] <= 0.799225607;
cosLookup[6726] <= 0.799167977;
cosLookup[6727] <= 0.799110339;
cosLookup[6728] <= 0.799052694;
cosLookup[6729] <= 0.798995042;
cosLookup[6730] <= 0.798937382;
cosLookup[6731] <= 0.798879715;
cosLookup[6732] <= 0.798822041;
cosLookup[6733] <= 0.798764359;
cosLookup[6734] <= 0.79870667;
cosLookup[6735] <= 0.798648974;
cosLookup[6736] <= 0.79859127;
cosLookup[6737] <= 0.798533559;
cosLookup[6738] <= 0.79847584;
cosLookup[6739] <= 0.798418114;
cosLookup[6740] <= 0.798360381;
cosLookup[6741] <= 0.798302641;
cosLookup[6742] <= 0.798244893;
cosLookup[6743] <= 0.798187138;
cosLookup[6744] <= 0.798129375;
cosLookup[6745] <= 0.798071606;
cosLookup[6746] <= 0.798013828;
cosLookup[6747] <= 0.797956044;
cosLookup[6748] <= 0.797898252;
cosLookup[6749] <= 0.797840453;
cosLookup[6750] <= 0.797782646;
cosLookup[6751] <= 0.797724833;
cosLookup[6752] <= 0.797667011;
cosLookup[6753] <= 0.797609183;
cosLookup[6754] <= 0.797551347;
cosLookup[6755] <= 0.797493504;
cosLookup[6756] <= 0.797435653;
cosLookup[6757] <= 0.797377796;
cosLookup[6758] <= 0.79731993;
cosLookup[6759] <= 0.797262058;
cosLookup[6760] <= 0.797204178;
cosLookup[6761] <= 0.797146291;
cosLookup[6762] <= 0.797088396;
cosLookup[6763] <= 0.797030495;
cosLookup[6764] <= 0.796972586;
cosLookup[6765] <= 0.796914669;
cosLookup[6766] <= 0.796856745;
cosLookup[6767] <= 0.796798814;
cosLookup[6768] <= 0.796740876;
cosLookup[6769] <= 0.79668293;
cosLookup[6770] <= 0.796624977;
cosLookup[6771] <= 0.796567017;
cosLookup[6772] <= 0.796509049;
cosLookup[6773] <= 0.796451074;
cosLookup[6774] <= 0.796393091;
cosLookup[6775] <= 0.796335102;
cosLookup[6776] <= 0.796277105;
cosLookup[6777] <= 0.7962191;
cosLookup[6778] <= 0.796161089;
cosLookup[6779] <= 0.79610307;
cosLookup[6780] <= 0.796045043;
cosLookup[6781] <= 0.79598701;
cosLookup[6782] <= 0.795928969;
cosLookup[6783] <= 0.795870921;
cosLookup[6784] <= 0.795812865;
cosLookup[6785] <= 0.795754802;
cosLookup[6786] <= 0.795696732;
cosLookup[6787] <= 0.795638655;
cosLookup[6788] <= 0.79558057;
cosLookup[6789] <= 0.795522478;
cosLookup[6790] <= 0.795464378;
cosLookup[6791] <= 0.795406271;
cosLookup[6792] <= 0.795348157;
cosLookup[6793] <= 0.795290036;
cosLookup[6794] <= 0.795231907;
cosLookup[6795] <= 0.795173771;
cosLookup[6796] <= 0.795115628;
cosLookup[6797] <= 0.795057477;
cosLookup[6798] <= 0.794999319;
cosLookup[6799] <= 0.794941154;
cosLookup[6800] <= 0.794882982;
cosLookup[6801] <= 0.794824802;
cosLookup[6802] <= 0.794766615;
cosLookup[6803] <= 0.79470842;
cosLookup[6804] <= 0.794650218;
cosLookup[6805] <= 0.794592009;
cosLookup[6806] <= 0.794533793;
cosLookup[6807] <= 0.794475569;
cosLookup[6808] <= 0.794417338;
cosLookup[6809] <= 0.7943591;
cosLookup[6810] <= 0.794300854;
cosLookup[6811] <= 0.794242601;
cosLookup[6812] <= 0.794184341;
cosLookup[6813] <= 0.794126074;
cosLookup[6814] <= 0.794067799;
cosLookup[6815] <= 0.794009517;
cosLookup[6816] <= 0.793951227;
cosLookup[6817] <= 0.793892931;
cosLookup[6818] <= 0.793834627;
cosLookup[6819] <= 0.793776315;
cosLookup[6820] <= 0.793717997;
cosLookup[6821] <= 0.793659671;
cosLookup[6822] <= 0.793601338;
cosLookup[6823] <= 0.793542997;
cosLookup[6824] <= 0.793484649;
cosLookup[6825] <= 0.793426294;
cosLookup[6826] <= 0.793367932;
cosLookup[6827] <= 0.793309562;
cosLookup[6828] <= 0.793251185;
cosLookup[6829] <= 0.793192801;
cosLookup[6830] <= 0.79313441;
cosLookup[6831] <= 0.793076011;
cosLookup[6832] <= 0.793017605;
cosLookup[6833] <= 0.792959191;
cosLookup[6834] <= 0.792900771;
cosLookup[6835] <= 0.792842343;
cosLookup[6836] <= 0.792783907;
cosLookup[6837] <= 0.792725465;
cosLookup[6838] <= 0.792667015;
cosLookup[6839] <= 0.792608558;
cosLookup[6840] <= 0.792550093;
cosLookup[6841] <= 0.792491622;
cosLookup[6842] <= 0.792433143;
cosLookup[6843] <= 0.792374656;
cosLookup[6844] <= 0.792316163;
cosLookup[6845] <= 0.792257662;
cosLookup[6846] <= 0.792199154;
cosLookup[6847] <= 0.792140638;
cosLookup[6848] <= 0.792082116;
cosLookup[6849] <= 0.792023586;
cosLookup[6850] <= 0.791965049;
cosLookup[6851] <= 0.791906504;
cosLookup[6852] <= 0.791847952;
cosLookup[6853] <= 0.791789393;
cosLookup[6854] <= 0.791730827;
cosLookup[6855] <= 0.791672253;
cosLookup[6856] <= 0.791613672;
cosLookup[6857] <= 0.791555084;
cosLookup[6858] <= 0.791496488;
cosLookup[6859] <= 0.791437886;
cosLookup[6860] <= 0.791379276;
cosLookup[6861] <= 0.791320658;
cosLookup[6862] <= 0.791262034;
cosLookup[6863] <= 0.791203402;
cosLookup[6864] <= 0.791144763;
cosLookup[6865] <= 0.791086116;
cosLookup[6866] <= 0.791027463;
cosLookup[6867] <= 0.790968802;
cosLookup[6868] <= 0.790910133;
cosLookup[6869] <= 0.790851458;
cosLookup[6870] <= 0.790792775;
cosLookup[6871] <= 0.790734085;
cosLookup[6872] <= 0.790675388;
cosLookup[6873] <= 0.790616683;
cosLookup[6874] <= 0.790557971;
cosLookup[6875] <= 0.790499252;
cosLookup[6876] <= 0.790440526;
cosLookup[6877] <= 0.790381792;
cosLookup[6878] <= 0.790323051;
cosLookup[6879] <= 0.790264303;
cosLookup[6880] <= 0.790205548;
cosLookup[6881] <= 0.790146785;
cosLookup[6882] <= 0.790088015;
cosLookup[6883] <= 0.790029238;
cosLookup[6884] <= 0.789970453;
cosLookup[6885] <= 0.789911662;
cosLookup[6886] <= 0.789852863;
cosLookup[6887] <= 0.789794056;
cosLookup[6888] <= 0.789735243;
cosLookup[6889] <= 0.789676422;
cosLookup[6890] <= 0.789617594;
cosLookup[6891] <= 0.789558759;
cosLookup[6892] <= 0.789499916;
cosLookup[6893] <= 0.789441066;
cosLookup[6894] <= 0.789382209;
cosLookup[6895] <= 0.789323345;
cosLookup[6896] <= 0.789264473;
cosLookup[6897] <= 0.789205594;
cosLookup[6898] <= 0.789146708;
cosLookup[6899] <= 0.789087815;
cosLookup[6900] <= 0.789028914;
cosLookup[6901] <= 0.788970007;
cosLookup[6902] <= 0.788911091;
cosLookup[6903] <= 0.788852169;
cosLookup[6904] <= 0.788793239;
cosLookup[6905] <= 0.788734302;
cosLookup[6906] <= 0.788675358;
cosLookup[6907] <= 0.788616407;
cosLookup[6908] <= 0.788557448;
cosLookup[6909] <= 0.788498482;
cosLookup[6910] <= 0.788439509;
cosLookup[6911] <= 0.788380529;
cosLookup[6912] <= 0.788321541;
cosLookup[6913] <= 0.788262546;
cosLookup[6914] <= 0.788203544;
cosLookup[6915] <= 0.788144535;
cosLookup[6916] <= 0.788085518;
cosLookup[6917] <= 0.788026495;
cosLookup[6918] <= 0.787967463;
cosLookup[6919] <= 0.787908425;
cosLookup[6920] <= 0.78784938;
cosLookup[6921] <= 0.787790327;
cosLookup[6922] <= 0.787731267;
cosLookup[6923] <= 0.787672199;
cosLookup[6924] <= 0.787613125;
cosLookup[6925] <= 0.787554043;
cosLookup[6926] <= 0.787494954;
cosLookup[6927] <= 0.787435858;
cosLookup[6928] <= 0.787376754;
cosLookup[6929] <= 0.787317643;
cosLookup[6930] <= 0.787258525;
cosLookup[6931] <= 0.7871994;
cosLookup[6932] <= 0.787140268;
cosLookup[6933] <= 0.787081128;
cosLookup[6934] <= 0.787021981;
cosLookup[6935] <= 0.786962827;
cosLookup[6936] <= 0.786903666;
cosLookup[6937] <= 0.786844497;
cosLookup[6938] <= 0.786785321;
cosLookup[6939] <= 0.786726138;
cosLookup[6940] <= 0.786666948;
cosLookup[6941] <= 0.78660775;
cosLookup[6942] <= 0.786548545;
cosLookup[6943] <= 0.786489333;
cosLookup[6944] <= 0.786430114;
cosLookup[6945] <= 0.786370887;
cosLookup[6946] <= 0.786311654;
cosLookup[6947] <= 0.786252413;
cosLookup[6948] <= 0.786193165;
cosLookup[6949] <= 0.786133909;
cosLookup[6950] <= 0.786074647;
cosLookup[6951] <= 0.786015377;
cosLookup[6952] <= 0.7859561;
cosLookup[6953] <= 0.785896815;
cosLookup[6954] <= 0.785837524;
cosLookup[6955] <= 0.785778225;
cosLookup[6956] <= 0.785718919;
cosLookup[6957] <= 0.785659606;
cosLookup[6958] <= 0.785600285;
cosLookup[6959] <= 0.785540958;
cosLookup[6960] <= 0.785481623;
cosLookup[6961] <= 0.785422281;
cosLookup[6962] <= 0.785362932;
cosLookup[6963] <= 0.785303575;
cosLookup[6964] <= 0.785244211;
cosLookup[6965] <= 0.78518484;
cosLookup[6966] <= 0.785125462;
cosLookup[6967] <= 0.785066077;
cosLookup[6968] <= 0.785006684;
cosLookup[6969] <= 0.784947284;
cosLookup[6970] <= 0.784887877;
cosLookup[6971] <= 0.784828463;
cosLookup[6972] <= 0.784769041;
cosLookup[6973] <= 0.784709613;
cosLookup[6974] <= 0.784650177;
cosLookup[6975] <= 0.784590734;
cosLookup[6976] <= 0.784531283;
cosLookup[6977] <= 0.784471826;
cosLookup[6978] <= 0.784412361;
cosLookup[6979] <= 0.784352889;
cosLookup[6980] <= 0.78429341;
cosLookup[6981] <= 0.784233924;
cosLookup[6982] <= 0.78417443;
cosLookup[6983] <= 0.784114929;
cosLookup[6984] <= 0.784055421;
cosLookup[6985] <= 0.783995906;
cosLookup[6986] <= 0.783936384;
cosLookup[6987] <= 0.783876854;
cosLookup[6988] <= 0.783817317;
cosLookup[6989] <= 0.783757773;
cosLookup[6990] <= 0.783698222;
cosLookup[6991] <= 0.783638663;
cosLookup[6992] <= 0.783579098;
cosLookup[6993] <= 0.783519525;
cosLookup[6994] <= 0.783459945;
cosLookup[6995] <= 0.783400357;
cosLookup[6996] <= 0.783340763;
cosLookup[6997] <= 0.783281161;
cosLookup[6998] <= 0.783221552;
cosLookup[6999] <= 0.783161936;
cosLookup[7000] <= 0.783102313;
cosLookup[7001] <= 0.783042683;
cosLookup[7002] <= 0.782983045;
cosLookup[7003] <= 0.7829234;
cosLookup[7004] <= 0.782863748;
cosLookup[7005] <= 0.782804089;
cosLookup[7006] <= 0.782744422;
cosLookup[7007] <= 0.782684749;
cosLookup[7008] <= 0.782625068;
cosLookup[7009] <= 0.78256538;
cosLookup[7010] <= 0.782505684;
cosLookup[7011] <= 0.782445982;
cosLookup[7012] <= 0.782386272;
cosLookup[7013] <= 0.782326556;
cosLookup[7014] <= 0.782266832;
cosLookup[7015] <= 0.7822071;
cosLookup[7016] <= 0.782147362;
cosLookup[7017] <= 0.782087616;
cosLookup[7018] <= 0.782027864;
cosLookup[7019] <= 0.781968104;
cosLookup[7020] <= 0.781908337;
cosLookup[7021] <= 0.781848562;
cosLookup[7022] <= 0.781788781;
cosLookup[7023] <= 0.781728992;
cosLookup[7024] <= 0.781669196;
cosLookup[7025] <= 0.781609393;
cosLookup[7026] <= 0.781549583;
cosLookup[7027] <= 0.781489765;
cosLookup[7028] <= 0.781429941;
cosLookup[7029] <= 0.781370109;
cosLookup[7030] <= 0.78131027;
cosLookup[7031] <= 0.781250424;
cosLookup[7032] <= 0.78119057;
cosLookup[7033] <= 0.78113071;
cosLookup[7034] <= 0.781070842;
cosLookup[7035] <= 0.781010967;
cosLookup[7036] <= 0.780951085;
cosLookup[7037] <= 0.780891196;
cosLookup[7038] <= 0.780831299;
cosLookup[7039] <= 0.780771396;
cosLookup[7040] <= 0.780711485;
cosLookup[7041] <= 0.780651567;
cosLookup[7042] <= 0.780591642;
cosLookup[7043] <= 0.780531709;
cosLookup[7044] <= 0.78047177;
cosLookup[7045] <= 0.780411823;
cosLookup[7046] <= 0.780351869;
cosLookup[7047] <= 0.780291908;
cosLookup[7048] <= 0.78023194;
cosLookup[7049] <= 0.780171965;
cosLookup[7050] <= 0.780111982;
cosLookup[7051] <= 0.780051992;
cosLookup[7052] <= 0.779991995;
cosLookup[7053] <= 0.779931991;
cosLookup[7054] <= 0.77987198;
cosLookup[7055] <= 0.779811962;
cosLookup[7056] <= 0.779751936;
cosLookup[7057] <= 0.779691903;
cosLookup[7058] <= 0.779631864;
cosLookup[7059] <= 0.779571816;
cosLookup[7060] <= 0.779511762;
cosLookup[7061] <= 0.779451701;
cosLookup[7062] <= 0.779391632;
cosLookup[7063] <= 0.779331557;
cosLookup[7064] <= 0.779271474;
cosLookup[7065] <= 0.779211384;
cosLookup[7066] <= 0.779151286;
cosLookup[7067] <= 0.779091182;
cosLookup[7068] <= 0.77903107;
cosLookup[7069] <= 0.778970952;
cosLookup[7070] <= 0.778910826;
cosLookup[7071] <= 0.778850693;
cosLookup[7072] <= 0.778790553;
cosLookup[7073] <= 0.778730405;
cosLookup[7074] <= 0.778670251;
cosLookup[7075] <= 0.778610089;
cosLookup[7076] <= 0.77854992;
cosLookup[7077] <= 0.778489744;
cosLookup[7078] <= 0.778429561;
cosLookup[7079] <= 0.778369371;
cosLookup[7080] <= 0.778309173;
cosLookup[7081] <= 0.778248969;
cosLookup[7082] <= 0.778188757;
cosLookup[7083] <= 0.778128538;
cosLookup[7084] <= 0.778068312;
cosLookup[7085] <= 0.778008079;
cosLookup[7086] <= 0.777947838;
cosLookup[7087] <= 0.777887591;
cosLookup[7088] <= 0.777827336;
cosLookup[7089] <= 0.777767074;
cosLookup[7090] <= 0.777706805;
cosLookup[7091] <= 0.777646529;
cosLookup[7092] <= 0.777586246;
cosLookup[7093] <= 0.777525955;
cosLookup[7094] <= 0.777465658;
cosLookup[7095] <= 0.777405353;
cosLookup[7096] <= 0.777345041;
cosLookup[7097] <= 0.777284722;
cosLookup[7098] <= 0.777224396;
cosLookup[7099] <= 0.777164063;
cosLookup[7100] <= 0.777103722;
cosLookup[7101] <= 0.777043375;
cosLookup[7102] <= 0.77698302;
cosLookup[7103] <= 0.776922658;
cosLookup[7104] <= 0.776862289;
cosLookup[7105] <= 0.776801913;
cosLookup[7106] <= 0.77674153;
cosLookup[7107] <= 0.776681139;
cosLookup[7108] <= 0.776620742;
cosLookup[7109] <= 0.776560337;
cosLookup[7110] <= 0.776499925;
cosLookup[7111] <= 0.776439506;
cosLookup[7112] <= 0.77637908;
cosLookup[7113] <= 0.776318647;
cosLookup[7114] <= 0.776258206;
cosLookup[7115] <= 0.776197759;
cosLookup[7116] <= 0.776137304;
cosLookup[7117] <= 0.776076842;
cosLookup[7118] <= 0.776016373;
cosLookup[7119] <= 0.775955897;
cosLookup[7120] <= 0.775895414;
cosLookup[7121] <= 0.775834924;
cosLookup[7122] <= 0.775774426;
cosLookup[7123] <= 0.775713922;
cosLookup[7124] <= 0.77565341;
cosLookup[7125] <= 0.775592891;
cosLookup[7126] <= 0.775532365;
cosLookup[7127] <= 0.775471832;
cosLookup[7128] <= 0.775411291;
cosLookup[7129] <= 0.775350744;
cosLookup[7130] <= 0.77529019;
cosLookup[7131] <= 0.775229628;
cosLookup[7132] <= 0.775169059;
cosLookup[7133] <= 0.775108483;
cosLookup[7134] <= 0.7750479;
cosLookup[7135] <= 0.77498731;
cosLookup[7136] <= 0.774926713;
cosLookup[7137] <= 0.774866108;
cosLookup[7138] <= 0.774805497;
cosLookup[7139] <= 0.774744878;
cosLookup[7140] <= 0.774684252;
cosLookup[7141] <= 0.77462362;
cosLookup[7142] <= 0.77456298;
cosLookup[7143] <= 0.774502332;
cosLookup[7144] <= 0.774441678;
cosLookup[7145] <= 0.774381017;
cosLookup[7146] <= 0.774320348;
cosLookup[7147] <= 0.774259673;
cosLookup[7148] <= 0.77419899;
cosLookup[7149] <= 0.7741383;
cosLookup[7150] <= 0.774077603;
cosLookup[7151] <= 0.774016899;
cosLookup[7152] <= 0.773956188;
cosLookup[7153] <= 0.77389547;
cosLookup[7154] <= 0.773834744;
cosLookup[7155] <= 0.773774012;
cosLookup[7156] <= 0.773713272;
cosLookup[7157] <= 0.773652525;
cosLookup[7158] <= 0.773591771;
cosLookup[7159] <= 0.77353101;
cosLookup[7160] <= 0.773470242;
cosLookup[7161] <= 0.773409467;
cosLookup[7162] <= 0.773348685;
cosLookup[7163] <= 0.773287895;
cosLookup[7164] <= 0.773227099;
cosLookup[7165] <= 0.773166295;
cosLookup[7166] <= 0.773105484;
cosLookup[7167] <= 0.773044667;
cosLookup[7168] <= 0.772983842;
cosLookup[7169] <= 0.772923009;
cosLookup[7170] <= 0.77286217;
cosLookup[7171] <= 0.772801324;
cosLookup[7172] <= 0.772740471;
cosLookup[7173] <= 0.77267961;
cosLookup[7174] <= 0.772618743;
cosLookup[7175] <= 0.772557868;
cosLookup[7176] <= 0.772496986;
cosLookup[7177] <= 0.772436097;
cosLookup[7178] <= 0.772375201;
cosLookup[7179] <= 0.772314298;
cosLookup[7180] <= 0.772253388;
cosLookup[7181] <= 0.772192471;
cosLookup[7182] <= 0.772131546;
cosLookup[7183] <= 0.772070615;
cosLookup[7184] <= 0.772009676;
cosLookup[7185] <= 0.77194873;
cosLookup[7186] <= 0.771887778;
cosLookup[7187] <= 0.771826818;
cosLookup[7188] <= 0.771765851;
cosLookup[7189] <= 0.771704877;
cosLookup[7190] <= 0.771643896;
cosLookup[7191] <= 0.771582907;
cosLookup[7192] <= 0.771521912;
cosLookup[7193] <= 0.77146091;
cosLookup[7194] <= 0.7713999;
cosLookup[7195] <= 0.771338883;
cosLookup[7196] <= 0.77127786;
cosLookup[7197] <= 0.771216829;
cosLookup[7198] <= 0.771155791;
cosLookup[7199] <= 0.771094746;
cosLookup[7200] <= 0.771033694;
cosLookup[7201] <= 0.770972635;
cosLookup[7202] <= 0.770911568;
cosLookup[7203] <= 0.770850495;
cosLookup[7204] <= 0.770789415;
cosLookup[7205] <= 0.770728327;
cosLookup[7206] <= 0.770667233;
cosLookup[7207] <= 0.770606131;
cosLookup[7208] <= 0.770545022;
cosLookup[7209] <= 0.770483906;
cosLookup[7210] <= 0.770422783;
cosLookup[7211] <= 0.770361653;
cosLookup[7212] <= 0.770300516;
cosLookup[7213] <= 0.770239372;
cosLookup[7214] <= 0.770178221;
cosLookup[7215] <= 0.770117062;
cosLookup[7216] <= 0.770055897;
cosLookup[7217] <= 0.769994725;
cosLookup[7218] <= 0.769933545;
cosLookup[7219] <= 0.769872358;
cosLookup[7220] <= 0.769811165;
cosLookup[7221] <= 0.769749964;
cosLookup[7222] <= 0.769688756;
cosLookup[7223] <= 0.769627541;
cosLookup[7224] <= 0.769566319;
cosLookup[7225] <= 0.76950509;
cosLookup[7226] <= 0.769443854;
cosLookup[7227] <= 0.76938261;
cosLookup[7228] <= 0.76932136;
cosLookup[7229] <= 0.769260103;
cosLookup[7230] <= 0.769198838;
cosLookup[7231] <= 0.769137567;
cosLookup[7232] <= 0.769076288;
cosLookup[7233] <= 0.769015002;
cosLookup[7234] <= 0.76895371;
cosLookup[7235] <= 0.76889241;
cosLookup[7236] <= 0.768831103;
cosLookup[7237] <= 0.768769789;
cosLookup[7238] <= 0.768708468;
cosLookup[7239] <= 0.76864714;
cosLookup[7240] <= 0.768585805;
cosLookup[7241] <= 0.768524462;
cosLookup[7242] <= 0.768463113;
cosLookup[7243] <= 0.768401757;
cosLookup[7244] <= 0.768340393;
cosLookup[7245] <= 0.768279023;
cosLookup[7246] <= 0.768217645;
cosLookup[7247] <= 0.768156261;
cosLookup[7248] <= 0.768094869;
cosLookup[7249] <= 0.76803347;
cosLookup[7250] <= 0.767972065;
cosLookup[7251] <= 0.767910652;
cosLookup[7252] <= 0.767849232;
cosLookup[7253] <= 0.767787805;
cosLookup[7254] <= 0.767726371;
cosLookup[7255] <= 0.76766493;
cosLookup[7256] <= 0.767603482;
cosLookup[7257] <= 0.767542026;
cosLookup[7258] <= 0.767480564;
cosLookup[7259] <= 0.767419095;
cosLookup[7260] <= 0.767357618;
cosLookup[7261] <= 0.767296135;
cosLookup[7262] <= 0.767234645;
cosLookup[7263] <= 0.767173147;
cosLookup[7264] <= 0.767111642;
cosLookup[7265] <= 0.767050131;
cosLookup[7266] <= 0.766988612;
cosLookup[7267] <= 0.766927086;
cosLookup[7268] <= 0.766865554;
cosLookup[7269] <= 0.766804014;
cosLookup[7270] <= 0.766742467;
cosLookup[7271] <= 0.766680913;
cosLookup[7272] <= 0.766619352;
cosLookup[7273] <= 0.766557784;
cosLookup[7274] <= 0.766496209;
cosLookup[7275] <= 0.766434627;
cosLookup[7276] <= 0.766373038;
cosLookup[7277] <= 0.766311441;
cosLookup[7278] <= 0.766249838;
cosLookup[7279] <= 0.766188228;
cosLookup[7280] <= 0.766126611;
cosLookup[7281] <= 0.766064986;
cosLookup[7282] <= 0.766003355;
cosLookup[7283] <= 0.765941716;
cosLookup[7284] <= 0.765880071;
cosLookup[7285] <= 0.765818418;
cosLookup[7286] <= 0.765756759;
cosLookup[7287] <= 0.765695092;
cosLookup[7288] <= 0.765633418;
cosLookup[7289] <= 0.765571738;
cosLookup[7290] <= 0.76551005;
cosLookup[7291] <= 0.765448355;
cosLookup[7292] <= 0.765386653;
cosLookup[7293] <= 0.765324944;
cosLookup[7294] <= 0.765263229;
cosLookup[7295] <= 0.765201506;
cosLookup[7296] <= 0.765139776;
cosLookup[7297] <= 0.765078039;
cosLookup[7298] <= 0.765016295;
cosLookup[7299] <= 0.764954544;
cosLookup[7300] <= 0.764892785;
cosLookup[7301] <= 0.76483102;
cosLookup[7302] <= 0.764769248;
cosLookup[7303] <= 0.764707469;
cosLookup[7304] <= 0.764645683;
cosLookup[7305] <= 0.76458389;
cosLookup[7306] <= 0.764522089;
cosLookup[7307] <= 0.764460282;
cosLookup[7308] <= 0.764398468;
cosLookup[7309] <= 0.764336646;
cosLookup[7310] <= 0.764274818;
cosLookup[7311] <= 0.764212982;
cosLookup[7312] <= 0.76415114;
cosLookup[7313] <= 0.764089291;
cosLookup[7314] <= 0.764027434;
cosLookup[7315] <= 0.763965571;
cosLookup[7316] <= 0.7639037;
cosLookup[7317] <= 0.763841823;
cosLookup[7318] <= 0.763779938;
cosLookup[7319] <= 0.763718046;
cosLookup[7320] <= 0.763656148;
cosLookup[7321] <= 0.763594242;
cosLookup[7322] <= 0.763532329;
cosLookup[7323] <= 0.76347041;
cosLookup[7324] <= 0.763408483;
cosLookup[7325] <= 0.763346549;
cosLookup[7326] <= 0.763284609;
cosLookup[7327] <= 0.763222661;
cosLookup[7328] <= 0.763160706;
cosLookup[7329] <= 0.763098744;
cosLookup[7330] <= 0.763036776;
cosLookup[7331] <= 0.7629748;
cosLookup[7332] <= 0.762912817;
cosLookup[7333] <= 0.762850827;
cosLookup[7334] <= 0.76278883;
cosLookup[7335] <= 0.762726826;
cosLookup[7336] <= 0.762664816;
cosLookup[7337] <= 0.762602798;
cosLookup[7338] <= 0.762540773;
cosLookup[7339] <= 0.762478741;
cosLookup[7340] <= 0.762416702;
cosLookup[7341] <= 0.762354656;
cosLookup[7342] <= 0.762292603;
cosLookup[7343] <= 0.762230543;
cosLookup[7344] <= 0.762168476;
cosLookup[7345] <= 0.762106402;
cosLookup[7346] <= 0.762044321;
cosLookup[7347] <= 0.761982233;
cosLookup[7348] <= 0.761920138;
cosLookup[7349] <= 0.761858036;
cosLookup[7350] <= 0.761795927;
cosLookup[7351] <= 0.761733811;
cosLookup[7352] <= 0.761671689;
cosLookup[7353] <= 0.761609559;
cosLookup[7354] <= 0.761547422;
cosLookup[7355] <= 0.761485278;
cosLookup[7356] <= 0.761423127;
cosLookup[7357] <= 0.761360969;
cosLookup[7358] <= 0.761298804;
cosLookup[7359] <= 0.761236632;
cosLookup[7360] <= 0.761174453;
cosLookup[7361] <= 0.761112267;
cosLookup[7362] <= 0.761050074;
cosLookup[7363] <= 0.760987874;
cosLookup[7364] <= 0.760925667;
cosLookup[7365] <= 0.760863453;
cosLookup[7366] <= 0.760801232;
cosLookup[7367] <= 0.760739004;
cosLookup[7368] <= 0.760676769;
cosLookup[7369] <= 0.760614527;
cosLookup[7370] <= 0.760552278;
cosLookup[7371] <= 0.760490022;
cosLookup[7372] <= 0.760427759;
cosLookup[7373] <= 0.760365489;
cosLookup[7374] <= 0.760303212;
cosLookup[7375] <= 0.760240929;
cosLookup[7376] <= 0.760178638;
cosLookup[7377] <= 0.76011634;
cosLookup[7378] <= 0.760054035;
cosLookup[7379] <= 0.759991723;
cosLookup[7380] <= 0.759929404;
cosLookup[7381] <= 0.759867079;
cosLookup[7382] <= 0.759804746;
cosLookup[7383] <= 0.759742406;
cosLookup[7384] <= 0.759680059;
cosLookup[7385] <= 0.759617706;
cosLookup[7386] <= 0.759555345;
cosLookup[7387] <= 0.759492977;
cosLookup[7388] <= 0.759430602;
cosLookup[7389] <= 0.759368221;
cosLookup[7390] <= 0.759305832;
cosLookup[7391] <= 0.759243436;
cosLookup[7392] <= 0.759181034;
cosLookup[7393] <= 0.759118624;
cosLookup[7394] <= 0.759056208;
cosLookup[7395] <= 0.758993784;
cosLookup[7396] <= 0.758931354;
cosLookup[7397] <= 0.758868916;
cosLookup[7398] <= 0.758806472;
cosLookup[7399] <= 0.75874402;
cosLookup[7400] <= 0.758681562;
cosLookup[7401] <= 0.758619096;
cosLookup[7402] <= 0.758556624;
cosLookup[7403] <= 0.758494145;
cosLookup[7404] <= 0.758431658;
cosLookup[7405] <= 0.758369165;
cosLookup[7406] <= 0.758306665;
cosLookup[7407] <= 0.758244157;
cosLookup[7408] <= 0.758181643;
cosLookup[7409] <= 0.758119122;
cosLookup[7410] <= 0.758056594;
cosLookup[7411] <= 0.757994059;
cosLookup[7412] <= 0.757931517;
cosLookup[7413] <= 0.757868968;
cosLookup[7414] <= 0.757806412;
cosLookup[7415] <= 0.757743849;
cosLookup[7416] <= 0.757681279;
cosLookup[7417] <= 0.757618702;
cosLookup[7418] <= 0.757556118;
cosLookup[7419] <= 0.757493527;
cosLookup[7420] <= 0.757430929;
cosLookup[7421] <= 0.757368324;
cosLookup[7422] <= 0.757305713;
cosLookup[7423] <= 0.757243094;
cosLookup[7424] <= 0.757180468;
cosLookup[7425] <= 0.757117836;
cosLookup[7426] <= 0.757055196;
cosLookup[7427] <= 0.75699255;
cosLookup[7428] <= 0.756929896;
cosLookup[7429] <= 0.756867236;
cosLookup[7430] <= 0.756804568;
cosLookup[7431] <= 0.756741894;
cosLookup[7432] <= 0.756679213;
cosLookup[7433] <= 0.756616524;
cosLookup[7434] <= 0.756553829;
cosLookup[7435] <= 0.756491127;
cosLookup[7436] <= 0.756428418;
cosLookup[7437] <= 0.756365702;
cosLookup[7438] <= 0.756302979;
cosLookup[7439] <= 0.756240249;
cosLookup[7440] <= 0.756177512;
cosLookup[7441] <= 0.756114768;
cosLookup[7442] <= 0.756052017;
cosLookup[7443] <= 0.755989259;
cosLookup[7444] <= 0.755926494;
cosLookup[7445] <= 0.755863723;
cosLookup[7446] <= 0.755800944;
cosLookup[7447] <= 0.755738158;
cosLookup[7448] <= 0.755675366;
cosLookup[7449] <= 0.755612566;
cosLookup[7450] <= 0.75554976;
cosLookup[7451] <= 0.755486946;
cosLookup[7452] <= 0.755424126;
cosLookup[7453] <= 0.755361299;
cosLookup[7454] <= 0.755298465;
cosLookup[7455] <= 0.755235623;
cosLookup[7456] <= 0.755172775;
cosLookup[7457] <= 0.75510992;
cosLookup[7458] <= 0.755047058;
cosLookup[7459] <= 0.754984189;
cosLookup[7460] <= 0.754921313;
cosLookup[7461] <= 0.754858431;
cosLookup[7462] <= 0.754795541;
cosLookup[7463] <= 0.754732644;
cosLookup[7464] <= 0.75466974;
cosLookup[7465] <= 0.75460683;
cosLookup[7466] <= 0.754543912;
cosLookup[7467] <= 0.754480988;
cosLookup[7468] <= 0.754418057;
cosLookup[7469] <= 0.754355118;
cosLookup[7470] <= 0.754292173;
cosLookup[7471] <= 0.754229221;
cosLookup[7472] <= 0.754166262;
cosLookup[7473] <= 0.754103296;
cosLookup[7474] <= 0.754040323;
cosLookup[7475] <= 0.753977343;
cosLookup[7476] <= 0.753914356;
cosLookup[7477] <= 0.753851362;
cosLookup[7478] <= 0.753788361;
cosLookup[7479] <= 0.753725354;
cosLookup[7480] <= 0.753662339;
cosLookup[7481] <= 0.753599318;
cosLookup[7482] <= 0.753536289;
cosLookup[7483] <= 0.753473254;
cosLookup[7484] <= 0.753410212;
cosLookup[7485] <= 0.753347162;
cosLookup[7486] <= 0.753284106;
cosLookup[7487] <= 0.753221043;
cosLookup[7488] <= 0.753157973;
cosLookup[7489] <= 0.753094896;
cosLookup[7490] <= 0.753031813;
cosLookup[7491] <= 0.752968722;
cosLookup[7492] <= 0.752905624;
cosLookup[7493] <= 0.752842519;
cosLookup[7494] <= 0.752779408;
cosLookup[7495] <= 0.75271629;
cosLookup[7496] <= 0.752653164;
cosLookup[7497] <= 0.752590032;
cosLookup[7498] <= 0.752526893;
cosLookup[7499] <= 0.752463747;
cosLookup[7500] <= 0.752400594;
cosLookup[7501] <= 0.752337434;
cosLookup[7502] <= 0.752274267;
cosLookup[7503] <= 0.752211093;
cosLookup[7504] <= 0.752147912;
cosLookup[7505] <= 0.752084725;
cosLookup[7506] <= 0.75202153;
cosLookup[7507] <= 0.751958329;
cosLookup[7508] <= 0.75189512;
cosLookup[7509] <= 0.751831905;
cosLookup[7510] <= 0.751768683;
cosLookup[7511] <= 0.751705454;
cosLookup[7512] <= 0.751642218;
cosLookup[7513] <= 0.751578975;
cosLookup[7514] <= 0.751515725;
cosLookup[7515] <= 0.751452469;
cosLookup[7516] <= 0.751389205;
cosLookup[7517] <= 0.751325934;
cosLookup[7518] <= 0.751262657;
cosLookup[7519] <= 0.751199373;
cosLookup[7520] <= 0.751136081;
cosLookup[7521] <= 0.751072783;
cosLookup[7522] <= 0.751009478;
cosLookup[7523] <= 0.750946166;
cosLookup[7524] <= 0.750882847;
cosLookup[7525] <= 0.750819522;
cosLookup[7526] <= 0.750756189;
cosLookup[7527] <= 0.750692849;
cosLookup[7528] <= 0.750629503;
cosLookup[7529] <= 0.750566149;
cosLookup[7530] <= 0.750502789;
cosLookup[7531] <= 0.750439422;
cosLookup[7532] <= 0.750376048;
cosLookup[7533] <= 0.750312667;
cosLookup[7534] <= 0.750249279;
cosLookup[7535] <= 0.750185884;
cosLookup[7536] <= 0.750122483;
cosLookup[7537] <= 0.750059074;
cosLookup[7538] <= 0.749995659;
cosLookup[7539] <= 0.749932236;
cosLookup[7540] <= 0.749868807;
cosLookup[7541] <= 0.749805371;
cosLookup[7542] <= 0.749741928;
cosLookup[7543] <= 0.749678478;
cosLookup[7544] <= 0.749615021;
cosLookup[7545] <= 0.749551557;
cosLookup[7546] <= 0.749488087;
cosLookup[7547] <= 0.749424609;
cosLookup[7548] <= 0.749361125;
cosLookup[7549] <= 0.749297634;
cosLookup[7550] <= 0.749234136;
cosLookup[7551] <= 0.749170631;
cosLookup[7552] <= 0.749107119;
cosLookup[7553] <= 0.7490436;
cosLookup[7554] <= 0.748980074;
cosLookup[7555] <= 0.748916542;
cosLookup[7556] <= 0.748853002;
cosLookup[7557] <= 0.748789456;
cosLookup[7558] <= 0.748725902;
cosLookup[7559] <= 0.748662342;
cosLookup[7560] <= 0.748598775;
cosLookup[7561] <= 0.748535201;
cosLookup[7562] <= 0.748471621;
cosLookup[7563] <= 0.748408033;
cosLookup[7564] <= 0.748344439;
cosLookup[7565] <= 0.748280837;
cosLookup[7566] <= 0.748217229;
cosLookup[7567] <= 0.748153614;
cosLookup[7568] <= 0.748089992;
cosLookup[7569] <= 0.748026363;
cosLookup[7570] <= 0.747962727;
cosLookup[7571] <= 0.747899084;
cosLookup[7572] <= 0.747835435;
cosLookup[7573] <= 0.747771778;
cosLookup[7574] <= 0.747708115;
cosLookup[7575] <= 0.747644445;
cosLookup[7576] <= 0.747580768;
cosLookup[7577] <= 0.747517084;
cosLookup[7578] <= 0.747453393;
cosLookup[7579] <= 0.747389696;
cosLookup[7580] <= 0.747325991;
cosLookup[7581] <= 0.74726228;
cosLookup[7582] <= 0.747198561;
cosLookup[7583] <= 0.747134836;
cosLookup[7584] <= 0.747071104;
cosLookup[7585] <= 0.747007365;
cosLookup[7586] <= 0.74694362;
cosLookup[7587] <= 0.746879867;
cosLookup[7588] <= 0.746816108;
cosLookup[7589] <= 0.746752341;
cosLookup[7590] <= 0.746688568;
cosLookup[7591] <= 0.746624788;
cosLookup[7592] <= 0.746561001;
cosLookup[7593] <= 0.746497207;
cosLookup[7594] <= 0.746433407;
cosLookup[7595] <= 0.746369599;
cosLookup[7596] <= 0.746305785;
cosLookup[7597] <= 0.746241963;
cosLookup[7598] <= 0.746178135;
cosLookup[7599] <= 0.7461143;
cosLookup[7600] <= 0.746050459;
cosLookup[7601] <= 0.74598661;
cosLookup[7602] <= 0.745922754;
cosLookup[7603] <= 0.745858892;
cosLookup[7604] <= 0.745795023;
cosLookup[7605] <= 0.745731147;
cosLookup[7606] <= 0.745667264;
cosLookup[7607] <= 0.745603374;
cosLookup[7608] <= 0.745539477;
cosLookup[7609] <= 0.745475574;
cosLookup[7610] <= 0.745411663;
cosLookup[7611] <= 0.745347746;
cosLookup[7612] <= 0.745283822;
cosLookup[7613] <= 0.745219891;
cosLookup[7614] <= 0.745155953;
cosLookup[7615] <= 0.745092009;
cosLookup[7616] <= 0.745028057;
cosLookup[7617] <= 0.744964099;
cosLookup[7618] <= 0.744900134;
cosLookup[7619] <= 0.744836162;
cosLookup[7620] <= 0.744772183;
cosLookup[7621] <= 0.744708197;
cosLookup[7622] <= 0.744644204;
cosLookup[7623] <= 0.744580205;
cosLookup[7624] <= 0.744516199;
cosLookup[7625] <= 0.744452186;
cosLookup[7626] <= 0.744388166;
cosLookup[7627] <= 0.744324139;
cosLookup[7628] <= 0.744260105;
cosLookup[7629] <= 0.744196065;
cosLookup[7630] <= 0.744132018;
cosLookup[7631] <= 0.744067963;
cosLookup[7632] <= 0.744003902;
cosLookup[7633] <= 0.743939835;
cosLookup[7634] <= 0.74387576;
cosLookup[7635] <= 0.743811678;
cosLookup[7636] <= 0.74374759;
cosLookup[7637] <= 0.743683495;
cosLookup[7638] <= 0.743619393;
cosLookup[7639] <= 0.743555284;
cosLookup[7640] <= 0.743491168;
cosLookup[7641] <= 0.743427046;
cosLookup[7642] <= 0.743362916;
cosLookup[7643] <= 0.74329878;
cosLookup[7644] <= 0.743234637;
cosLookup[7645] <= 0.743170487;
cosLookup[7646] <= 0.743106331;
cosLookup[7647] <= 0.743042167;
cosLookup[7648] <= 0.742977997;
cosLookup[7649] <= 0.74291382;
cosLookup[7650] <= 0.742849636;
cosLookup[7651] <= 0.742785445;
cosLookup[7652] <= 0.742721247;
cosLookup[7653] <= 0.742657043;
cosLookup[7654] <= 0.742592831;
cosLookup[7655] <= 0.742528613;
cosLookup[7656] <= 0.742464388;
cosLookup[7657] <= 0.742400156;
cosLookup[7658] <= 0.742335918;
cosLookup[7659] <= 0.742271672;
cosLookup[7660] <= 0.74220742;
cosLookup[7661] <= 0.742143161;
cosLookup[7662] <= 0.742078895;
cosLookup[7663] <= 0.742014622;
cosLookup[7664] <= 0.741950343;
cosLookup[7665] <= 0.741886056;
cosLookup[7666] <= 0.741821763;
cosLookup[7667] <= 0.741757463;
cosLookup[7668] <= 0.741693156;
cosLookup[7669] <= 0.741628842;
cosLookup[7670] <= 0.741564522;
cosLookup[7671] <= 0.741500195;
cosLookup[7672] <= 0.741435861;
cosLookup[7673] <= 0.74137152;
cosLookup[7674] <= 0.741307172;
cosLookup[7675] <= 0.741242817;
cosLookup[7676] <= 0.741178456;
cosLookup[7677] <= 0.741114088;
cosLookup[7678] <= 0.741049713;
cosLookup[7679] <= 0.740985331;
cosLookup[7680] <= 0.740920942;
cosLookup[7681] <= 0.740856547;
cosLookup[7682] <= 0.740792145;
cosLookup[7683] <= 0.740727736;
cosLookup[7684] <= 0.74066332;
cosLookup[7685] <= 0.740598897;
cosLookup[7686] <= 0.740534468;
cosLookup[7687] <= 0.740470031;
cosLookup[7688] <= 0.740405588;
cosLookup[7689] <= 0.740341138;
cosLookup[7690] <= 0.740276682;
cosLookup[7691] <= 0.740212218;
cosLookup[7692] <= 0.740147748;
cosLookup[7693] <= 0.740083271;
cosLookup[7694] <= 0.740018787;
cosLookup[7695] <= 0.739954296;
cosLookup[7696] <= 0.739889798;
cosLookup[7697] <= 0.739825294;
cosLookup[7698] <= 0.739760783;
cosLookup[7699] <= 0.739696265;
cosLookup[7700] <= 0.73963174;
cosLookup[7701] <= 0.739567209;
cosLookup[7702] <= 0.73950267;
cosLookup[7703] <= 0.739438125;
cosLookup[7704] <= 0.739373573;
cosLookup[7705] <= 0.739309015;
cosLookup[7706] <= 0.739244449;
cosLookup[7707] <= 0.739179877;
cosLookup[7708] <= 0.739115298;
cosLookup[7709] <= 0.739050712;
cosLookup[7710] <= 0.738986119;
cosLookup[7711] <= 0.73892152;
cosLookup[7712] <= 0.738856913;
cosLookup[7713] <= 0.7387923;
cosLookup[7714] <= 0.73872768;
cosLookup[7715] <= 0.738663054;
cosLookup[7716] <= 0.73859842;
cosLookup[7717] <= 0.73853378;
cosLookup[7718] <= 0.738469133;
cosLookup[7719] <= 0.738404479;
cosLookup[7720] <= 0.738339818;
cosLookup[7721] <= 0.738275151;
cosLookup[7722] <= 0.738210477;
cosLookup[7723] <= 0.738145796;
cosLookup[7724] <= 0.738081108;
cosLookup[7725] <= 0.738016414;
cosLookup[7726] <= 0.737951712;
cosLookup[7727] <= 0.737887004;
cosLookup[7728] <= 0.737822289;
cosLookup[7729] <= 0.737757568;
cosLookup[7730] <= 0.737692839;
cosLookup[7731] <= 0.737628104;
cosLookup[7732] <= 0.737563362;
cosLookup[7733] <= 0.737498613;
cosLookup[7734] <= 0.737433857;
cosLookup[7735] <= 0.737369095;
cosLookup[7736] <= 0.737304326;
cosLookup[7737] <= 0.73723955;
cosLookup[7738] <= 0.737174767;
cosLookup[7739] <= 0.737109978;
cosLookup[7740] <= 0.737045182;
cosLookup[7741] <= 0.736980379;
cosLookup[7742] <= 0.736915569;
cosLookup[7743] <= 0.736850752;
cosLookup[7744] <= 0.736785929;
cosLookup[7745] <= 0.736721099;
cosLookup[7746] <= 0.736656262;
cosLookup[7747] <= 0.736591418;
cosLookup[7748] <= 0.736526568;
cosLookup[7749] <= 0.736461711;
cosLookup[7750] <= 0.736396847;
cosLookup[7751] <= 0.736331976;
cosLookup[7752] <= 0.736267098;
cosLookup[7753] <= 0.736202214;
cosLookup[7754] <= 0.736137323;
cosLookup[7755] <= 0.736072425;
cosLookup[7756] <= 0.736007521;
cosLookup[7757] <= 0.735942609;
cosLookup[7758] <= 0.735877691;
cosLookup[7759] <= 0.735812766;
cosLookup[7760] <= 0.735747835;
cosLookup[7761] <= 0.735682896;
cosLookup[7762] <= 0.735617951;
cosLookup[7763] <= 0.735552999;
cosLookup[7764] <= 0.73548804;
cosLookup[7765] <= 0.735423075;
cosLookup[7766] <= 0.735358103;
cosLookup[7767] <= 0.735293124;
cosLookup[7768] <= 0.735228138;
cosLookup[7769] <= 0.735163145;
cosLookup[7770] <= 0.735098146;
cosLookup[7771] <= 0.73503314;
cosLookup[7772] <= 0.734968127;
cosLookup[7773] <= 0.734903108;
cosLookup[7774] <= 0.734838082;
cosLookup[7775] <= 0.734773049;
cosLookup[7776] <= 0.734708009;
cosLookup[7777] <= 0.734642962;
cosLookup[7778] <= 0.734577909;
cosLookup[7779] <= 0.734512849;
cosLookup[7780] <= 0.734447782;
cosLookup[7781] <= 0.734382708;
cosLookup[7782] <= 0.734317628;
cosLookup[7783] <= 0.734252541;
cosLookup[7784] <= 0.734187447;
cosLookup[7785] <= 0.734122347;
cosLookup[7786] <= 0.734057239;
cosLookup[7787] <= 0.733992125;
cosLookup[7788] <= 0.733927005;
cosLookup[7789] <= 0.733861877;
cosLookup[7790] <= 0.733796743;
cosLookup[7791] <= 0.733731602;
cosLookup[7792] <= 0.733666454;
cosLookup[7793] <= 0.733601299;
cosLookup[7794] <= 0.733536138;
cosLookup[7795] <= 0.73347097;
cosLookup[7796] <= 0.733405795;
cosLookup[7797] <= 0.733340614;
cosLookup[7798] <= 0.733275426;
cosLookup[7799] <= 0.733210231;
cosLookup[7800] <= 0.733145029;
cosLookup[7801] <= 0.73307982;
cosLookup[7802] <= 0.733014605;
cosLookup[7803] <= 0.732949383;
cosLookup[7804] <= 0.732884155;
cosLookup[7805] <= 0.732818919;
cosLookup[7806] <= 0.732753677;
cosLookup[7807] <= 0.732688428;
cosLookup[7808] <= 0.732623172;
cosLookup[7809] <= 0.73255791;
cosLookup[7810] <= 0.732492641;
cosLookup[7811] <= 0.732427365;
cosLookup[7812] <= 0.732362083;
cosLookup[7813] <= 0.732296793;
cosLookup[7814] <= 0.732231497;
cosLookup[7815] <= 0.732166195;
cosLookup[7816] <= 0.732100885;
cosLookup[7817] <= 0.732035569;
cosLookup[7818] <= 0.731970246;
cosLookup[7819] <= 0.731904916;
cosLookup[7820] <= 0.73183958;
cosLookup[7821] <= 0.731774237;
cosLookup[7822] <= 0.731708887;
cosLookup[7823] <= 0.73164353;
cosLookup[7824] <= 0.731578167;
cosLookup[7825] <= 0.731512797;
cosLookup[7826] <= 0.73144742;
cosLookup[7827] <= 0.731382037;
cosLookup[7828] <= 0.731316646;
cosLookup[7829] <= 0.731251249;
cosLookup[7830] <= 0.731185846;
cosLookup[7831] <= 0.731120435;
cosLookup[7832] <= 0.731055018;
cosLookup[7833] <= 0.730989594;
cosLookup[7834] <= 0.730924164;
cosLookup[7835] <= 0.730858727;
cosLookup[7836] <= 0.730793283;
cosLookup[7837] <= 0.730727832;
cosLookup[7838] <= 0.730662375;
cosLookup[7839] <= 0.73059691;
cosLookup[7840] <= 0.73053144;
cosLookup[7841] <= 0.730465962;
cosLookup[7842] <= 0.730400478;
cosLookup[7843] <= 0.730334987;
cosLookup[7844] <= 0.730269489;
cosLookup[7845] <= 0.730203985;
cosLookup[7846] <= 0.730138473;
cosLookup[7847] <= 0.730072956;
cosLookup[7848] <= 0.730007431;
cosLookup[7849] <= 0.7299419;
cosLookup[7850] <= 0.729876362;
cosLookup[7851] <= 0.729810817;
cosLookup[7852] <= 0.729745266;
cosLookup[7853] <= 0.729679708;
cosLookup[7854] <= 0.729614143;
cosLookup[7855] <= 0.729548571;
cosLookup[7856] <= 0.729482993;
cosLookup[7857] <= 0.729417408;
cosLookup[7858] <= 0.729351816;
cosLookup[7859] <= 0.729286218;
cosLookup[7860] <= 0.729220613;
cosLookup[7861] <= 0.729155001;
cosLookup[7862] <= 0.729089383;
cosLookup[7863] <= 0.729023758;
cosLookup[7864] <= 0.728958126;
cosLookup[7865] <= 0.728892487;
cosLookup[7866] <= 0.728826842;
cosLookup[7867] <= 0.72876119;
cosLookup[7868] <= 0.728695531;
cosLookup[7869] <= 0.728629866;
cosLookup[7870] <= 0.728564194;
cosLookup[7871] <= 0.728498515;
cosLookup[7872] <= 0.72843283;
cosLookup[7873] <= 0.728367138;
cosLookup[7874] <= 0.728301439;
cosLookup[7875] <= 0.728235733;
cosLookup[7876] <= 0.728170021;
cosLookup[7877] <= 0.728104302;
cosLookup[7878] <= 0.728038576;
cosLookup[7879] <= 0.727972844;
cosLookup[7880] <= 0.727907105;
cosLookup[7881] <= 0.727841359;
cosLookup[7882] <= 0.727775607;
cosLookup[7883] <= 0.727709848;
cosLookup[7884] <= 0.727644082;
cosLookup[7885] <= 0.72757831;
cosLookup[7886] <= 0.727512531;
cosLookup[7887] <= 0.727446745;
cosLookup[7888] <= 0.727380952;
cosLookup[7889] <= 0.727315153;
cosLookup[7890] <= 0.727249347;
cosLookup[7891] <= 0.727183535;
cosLookup[7892] <= 0.727117715;
cosLookup[7893] <= 0.727051889;
cosLookup[7894] <= 0.726986057;
cosLookup[7895] <= 0.726920217;
cosLookup[7896] <= 0.726854371;
cosLookup[7897] <= 0.726788519;
cosLookup[7898] <= 0.726722659;
cosLookup[7899] <= 0.726656793;
cosLookup[7900] <= 0.726590921;
cosLookup[7901] <= 0.726525041;
cosLookup[7902] <= 0.726459155;
cosLookup[7903] <= 0.726393262;
cosLookup[7904] <= 0.726327363;
cosLookup[7905] <= 0.726261457;
cosLookup[7906] <= 0.726195544;
cosLookup[7907] <= 0.726129625;
cosLookup[7908] <= 0.726063698;
cosLookup[7909] <= 0.725997766;
cosLookup[7910] <= 0.725931826;
cosLookup[7911] <= 0.72586588;
cosLookup[7912] <= 0.725799927;
cosLookup[7913] <= 0.725733968;
cosLookup[7914] <= 0.725668001;
cosLookup[7915] <= 0.725602029;
cosLookup[7916] <= 0.725536049;
cosLookup[7917] <= 0.725470063;
cosLookup[7918] <= 0.72540407;
cosLookup[7919] <= 0.72533807;
cosLookup[7920] <= 0.725272064;
cosLookup[7921] <= 0.725206051;
cosLookup[7922] <= 0.725140032;
cosLookup[7923] <= 0.725074006;
cosLookup[7924] <= 0.725007973;
cosLookup[7925] <= 0.724941933;
cosLookup[7926] <= 0.724875887;
cosLookup[7927] <= 0.724809834;
cosLookup[7928] <= 0.724743775;
cosLookup[7929] <= 0.724677709;
cosLookup[7930] <= 0.724611636;
cosLookup[7931] <= 0.724545556;
cosLookup[7932] <= 0.72447947;
cosLookup[7933] <= 0.724413377;
cosLookup[7934] <= 0.724347278;
cosLookup[7935] <= 0.724281172;
cosLookup[7936] <= 0.724215059;
cosLookup[7937] <= 0.724148939;
cosLookup[7938] <= 0.724082813;
cosLookup[7939] <= 0.72401668;
cosLookup[7940] <= 0.723950541;
cosLookup[7941] <= 0.723884395;
cosLookup[7942] <= 0.723818242;
cosLookup[7943] <= 0.723752083;
cosLookup[7944] <= 0.723685917;
cosLookup[7945] <= 0.723619744;
cosLookup[7946] <= 0.723553565;
cosLookup[7947] <= 0.723487379;
cosLookup[7948] <= 0.723421186;
cosLookup[7949] <= 0.723354987;
cosLookup[7950] <= 0.723288781;
cosLookup[7951] <= 0.723222568;
cosLookup[7952] <= 0.723156349;
cosLookup[7953] <= 0.723090123;
cosLookup[7954] <= 0.72302389;
cosLookup[7955] <= 0.722957651;
cosLookup[7956] <= 0.722891405;
cosLookup[7957] <= 0.722825153;
cosLookup[7958] <= 0.722758894;
cosLookup[7959] <= 0.722692628;
cosLookup[7960] <= 0.722626356;
cosLookup[7961] <= 0.722560077;
cosLookup[7962] <= 0.722493791;
cosLookup[7963] <= 0.722427498;
cosLookup[7964] <= 0.722361199;
cosLookup[7965] <= 0.722294894;
cosLookup[7966] <= 0.722228582;
cosLookup[7967] <= 0.722162263;
cosLookup[7968] <= 0.722095937;
cosLookup[7969] <= 0.722029605;
cosLookup[7970] <= 0.721963266;
cosLookup[7971] <= 0.721896921;
cosLookup[7972] <= 0.721830569;
cosLookup[7973] <= 0.72176421;
cosLookup[7974] <= 0.721697844;
cosLookup[7975] <= 0.721631472;
cosLookup[7976] <= 0.721565094;
cosLookup[7977] <= 0.721498709;
cosLookup[7978] <= 0.721432317;
cosLookup[7979] <= 0.721365918;
cosLookup[7980] <= 0.721299513;
cosLookup[7981] <= 0.721233101;
cosLookup[7982] <= 0.721166683;
cosLookup[7983] <= 0.721100258;
cosLookup[7984] <= 0.721033826;
cosLookup[7985] <= 0.720967388;
cosLookup[7986] <= 0.720900943;
cosLookup[7987] <= 0.720834491;
cosLookup[7988] <= 0.720768033;
cosLookup[7989] <= 0.720701568;
cosLookup[7990] <= 0.720635097;
cosLookup[7991] <= 0.720568619;
cosLookup[7992] <= 0.720502134;
cosLookup[7993] <= 0.720435643;
cosLookup[7994] <= 0.720369145;
cosLookup[7995] <= 0.72030264;
cosLookup[7996] <= 0.720236129;
cosLookup[7997] <= 0.720169611;
cosLookup[7998] <= 0.720103087;
cosLookup[7999] <= 0.720036556;
cosLookup[8000] <= 0.719970018;
cosLookup[8001] <= 0.719903474;
cosLookup[8002] <= 0.719836923;
cosLookup[8003] <= 0.719770365;
cosLookup[8004] <= 0.719703801;
cosLookup[8005] <= 0.71963723;
cosLookup[8006] <= 0.719570653;
cosLookup[8007] <= 0.719504069;
cosLookup[8008] <= 0.719437479;
cosLookup[8009] <= 0.719370881;
cosLookup[8010] <= 0.719304277;
cosLookup[8011] <= 0.719237667;
cosLookup[8012] <= 0.71917105;
cosLookup[8013] <= 0.719104426;
cosLookup[8014] <= 0.719037796;
cosLookup[8015] <= 0.718971159;
cosLookup[8016] <= 0.718904516;
cosLookup[8017] <= 0.718837866;
cosLookup[8018] <= 0.718771209;
cosLookup[8019] <= 0.718704546;
cosLookup[8020] <= 0.718637876;
cosLookup[8021] <= 0.718571199;
cosLookup[8022] <= 0.718504516;
cosLookup[8023] <= 0.718437826;
cosLookup[8024] <= 0.71837113;
cosLookup[8025] <= 0.718304427;
cosLookup[8026] <= 0.718237717;
cosLookup[8027] <= 0.718171001;
cosLookup[8028] <= 0.718104279;
cosLookup[8029] <= 0.718037549;
cosLookup[8030] <= 0.717970813;
cosLookup[8031] <= 0.717904071;
cosLookup[8032] <= 0.717837322;
cosLookup[8033] <= 0.717770566;
cosLookup[8034] <= 0.717703803;
cosLookup[8035] <= 0.717637034;
cosLookup[8036] <= 0.717570259;
cosLookup[8037] <= 0.717503477;
cosLookup[8038] <= 0.717436688;
cosLookup[8039] <= 0.717369893;
cosLookup[8040] <= 0.717303091;
cosLookup[8041] <= 0.717236282;
cosLookup[8042] <= 0.717169467;
cosLookup[8043] <= 0.717102645;
cosLookup[8044] <= 0.717035817;
cosLookup[8045] <= 0.716968982;
cosLookup[8046] <= 0.716902141;
cosLookup[8047] <= 0.716835293;
cosLookup[8048] <= 0.716768438;
cosLookup[8049] <= 0.716701577;
cosLookup[8050] <= 0.716634709;
cosLookup[8051] <= 0.716567834;
cosLookup[8052] <= 0.716500953;
cosLookup[8053] <= 0.716434066;
cosLookup[8054] <= 0.716367172;
cosLookup[8055] <= 0.716300271;
cosLookup[8056] <= 0.716233363;
cosLookup[8057] <= 0.71616645;
cosLookup[8058] <= 0.716099529;
cosLookup[8059] <= 0.716032602;
cosLookup[8060] <= 0.715965668;
cosLookup[8061] <= 0.715898728;
cosLookup[8062] <= 0.715831781;
cosLookup[8063] <= 0.715764828;
cosLookup[8064] <= 0.715697868;
cosLookup[8065] <= 0.715630901;
cosLookup[8066] <= 0.715563928;
cosLookup[8067] <= 0.715496948;
cosLookup[8068] <= 0.715429962;
cosLookup[8069] <= 0.715362969;
cosLookup[8070] <= 0.715295969;
cosLookup[8071] <= 0.715228963;
cosLookup[8072] <= 0.715161951;
cosLookup[8073] <= 0.715094931;
cosLookup[8074] <= 0.715027906;
cosLookup[8075] <= 0.714960873;
cosLookup[8076] <= 0.714893834;
cosLookup[8077] <= 0.714826789;
cosLookup[8078] <= 0.714759737;
cosLookup[8079] <= 0.714692678;
cosLookup[8080] <= 0.714625613;
cosLookup[8081] <= 0.714558541;
cosLookup[8082] <= 0.714491463;
cosLookup[8083] <= 0.714424378;
cosLookup[8084] <= 0.714357286;
cosLookup[8085] <= 0.714290188;
cosLookup[8086] <= 0.714223084;
cosLookup[8087] <= 0.714155972;
cosLookup[8088] <= 0.714088855;
cosLookup[8089] <= 0.71402173;
cosLookup[8090] <= 0.7139546;
cosLookup[8091] <= 0.713887462;
cosLookup[8092] <= 0.713820318;
cosLookup[8093] <= 0.713753167;
cosLookup[8094] <= 0.71368601;
cosLookup[8095] <= 0.713618847;
cosLookup[8096] <= 0.713551676;
cosLookup[8097] <= 0.7134845;
cosLookup[8098] <= 0.713417316;
cosLookup[8099] <= 0.713350126;
cosLookup[8100] <= 0.71328293;
cosLookup[8101] <= 0.713215727;
cosLookup[8102] <= 0.713148517;
cosLookup[8103] <= 0.713081301;
cosLookup[8104] <= 0.713014078;
cosLookup[8105] <= 0.712946849;
cosLookup[8106] <= 0.712879613;
cosLookup[8107] <= 0.712812371;
cosLookup[8108] <= 0.712745122;
cosLookup[8109] <= 0.712677866;
cosLookup[8110] <= 0.712610604;
cosLookup[8111] <= 0.712543336;
cosLookup[8112] <= 0.712476061;
cosLookup[8113] <= 0.712408779;
cosLookup[8114] <= 0.712341491;
cosLookup[8115] <= 0.712274196;
cosLookup[8116] <= 0.712206895;
cosLookup[8117] <= 0.712139587;
cosLookup[8118] <= 0.712072272;
cosLookup[8119] <= 0.712004951;
cosLookup[8120] <= 0.711937624;
cosLookup[8121] <= 0.71187029;
cosLookup[8122] <= 0.711802949;
cosLookup[8123] <= 0.711735602;
cosLookup[8124] <= 0.711668248;
cosLookup[8125] <= 0.711600888;
cosLookup[8126] <= 0.711533521;
cosLookup[8127] <= 0.711466148;
cosLookup[8128] <= 0.711398768;
cosLookup[8129] <= 0.711331382;
cosLookup[8130] <= 0.711263989;
cosLookup[8131] <= 0.711196589;
cosLookup[8132] <= 0.711129183;
cosLookup[8133] <= 0.711061771;
cosLookup[8134] <= 0.710994352;
cosLookup[8135] <= 0.710926926;
cosLookup[8136] <= 0.710859494;
cosLookup[8137] <= 0.710792055;
cosLookup[8138] <= 0.71072461;
cosLookup[8139] <= 0.710657158;
cosLookup[8140] <= 0.7105897;
cosLookup[8141] <= 0.710522235;
cosLookup[8142] <= 0.710454764;
cosLookup[8143] <= 0.710387286;
cosLookup[8144] <= 0.710319802;
cosLookup[8145] <= 0.710252311;
cosLookup[8146] <= 0.710184813;
cosLookup[8147] <= 0.710117309;
cosLookup[8148] <= 0.710049799;
cosLookup[8149] <= 0.709982282;
cosLookup[8150] <= 0.709914758;
cosLookup[8151] <= 0.709847228;
cosLookup[8152] <= 0.709779691;
cosLookup[8153] <= 0.709712148;
cosLookup[8154] <= 0.709644598;
cosLookup[8155] <= 0.709577042;
cosLookup[8156] <= 0.709509479;
cosLookup[8157] <= 0.70944191;
cosLookup[8158] <= 0.709374334;
cosLookup[8159] <= 0.709306752;
cosLookup[8160] <= 0.709239163;
cosLookup[8161] <= 0.709171568;
cosLookup[8162] <= 0.709103966;
cosLookup[8163] <= 0.709036358;
cosLookup[8164] <= 0.708968743;
cosLookup[8165] <= 0.708901121;
cosLookup[8166] <= 0.708833493;
cosLookup[8167] <= 0.708765859;
cosLookup[8168] <= 0.708698218;
cosLookup[8169] <= 0.708630571;
cosLookup[8170] <= 0.708562917;
cosLookup[8171] <= 0.708495256;
cosLookup[8172] <= 0.708427589;
cosLookup[8173] <= 0.708359915;
cosLookup[8174] <= 0.708292235;
cosLookup[8175] <= 0.708224549;
cosLookup[8176] <= 0.708156856;
cosLookup[8177] <= 0.708089156;
cosLookup[8178] <= 0.70802145;
cosLookup[8179] <= 0.707953738;
cosLookup[8180] <= 0.707886018;
cosLookup[8181] <= 0.707818293;
cosLookup[8182] <= 0.707750561;
cosLookup[8183] <= 0.707682822;
cosLookup[8184] <= 0.707615077;
cosLookup[8185] <= 0.707547325;
cosLookup[8186] <= 0.707479567;
cosLookup[8187] <= 0.707411803;
cosLookup[8188] <= 0.707344031;
cosLookup[8189] <= 0.707276254;
cosLookup[8190] <= 0.70720847;
cosLookup[8191] <= 0.707140679;
cosLookup[8192] <= 0.707072882;
cosLookup[8193] <= 0.707005078;
cosLookup[8194] <= 0.706937268;
cosLookup[8195] <= 0.706869451;
cosLookup[8196] <= 0.706801628;
cosLookup[8197] <= 0.706733799;
cosLookup[8198] <= 0.706665962;
cosLookup[8199] <= 0.70659812;
cosLookup[8200] <= 0.706530271;
cosLookup[8201] <= 0.706462415;
cosLookup[8202] <= 0.706394553;
cosLookup[8203] <= 0.706326684;
cosLookup[8204] <= 0.706258809;
cosLookup[8205] <= 0.706190928;
cosLookup[8206] <= 0.706123039;
cosLookup[8207] <= 0.706055145;
cosLookup[8208] <= 0.705987244;
cosLookup[8209] <= 0.705919336;
cosLookup[8210] <= 0.705851422;
cosLookup[8211] <= 0.705783502;
cosLookup[8212] <= 0.705715575;
cosLookup[8213] <= 0.705647641;
cosLookup[8214] <= 0.705579701;
cosLookup[8215] <= 0.705511755;
cosLookup[8216] <= 0.705443802;
cosLookup[8217] <= 0.705375842;
cosLookup[8218] <= 0.705307876;
cosLookup[8219] <= 0.705239904;
cosLookup[8220] <= 0.705171925;
cosLookup[8221] <= 0.705103939;
cosLookup[8222] <= 0.705035948;
cosLookup[8223] <= 0.704967949;
cosLookup[8224] <= 0.704899944;
cosLookup[8225] <= 0.704831933;
cosLookup[8226] <= 0.704763915;
cosLookup[8227] <= 0.704695891;
cosLookup[8228] <= 0.70462786;
cosLookup[8229] <= 0.704559823;
cosLookup[8230] <= 0.704491779;
cosLookup[8231] <= 0.704423729;
cosLookup[8232] <= 0.704355672;
cosLookup[8233] <= 0.704287609;
cosLookup[8234] <= 0.70421954;
cosLookup[8235] <= 0.704151463;
cosLookup[8236] <= 0.704083381;
cosLookup[8237] <= 0.704015292;
cosLookup[8238] <= 0.703947196;
cosLookup[8239] <= 0.703879094;
cosLookup[8240] <= 0.703810986;
cosLookup[8241] <= 0.703742871;
cosLookup[8242] <= 0.70367475;
cosLookup[8243] <= 0.703606622;
cosLookup[8244] <= 0.703538487;
cosLookup[8245] <= 0.703470347;
cosLookup[8246] <= 0.703402199;
cosLookup[8247] <= 0.703334046;
cosLookup[8248] <= 0.703265885;
cosLookup[8249] <= 0.703197719;
cosLookup[8250] <= 0.703129546;
cosLookup[8251] <= 0.703061366;
cosLookup[8252] <= 0.70299318;
cosLookup[8253] <= 0.702924988;
cosLookup[8254] <= 0.702856789;
cosLookup[8255] <= 0.702788583;
cosLookup[8256] <= 0.702720371;
cosLookup[8257] <= 0.702652153;
cosLookup[8258] <= 0.702583928;
cosLookup[8259] <= 0.702515697;
cosLookup[8260] <= 0.702447459;
cosLookup[8261] <= 0.702379215;
cosLookup[8262] <= 0.702310964;
cosLookup[8263] <= 0.702242707;
cosLookup[8264] <= 0.702174444;
cosLookup[8265] <= 0.702106174;
cosLookup[8266] <= 0.702037897;
cosLookup[8267] <= 0.701969614;
cosLookup[8268] <= 0.701901325;
cosLookup[8269] <= 0.701833029;
cosLookup[8270] <= 0.701764727;
cosLookup[8271] <= 0.701696418;
cosLookup[8272] <= 0.701628103;
cosLookup[8273] <= 0.701559781;
cosLookup[8274] <= 0.701491453;
cosLookup[8275] <= 0.701423119;
cosLookup[8276] <= 0.701354778;
cosLookup[8277] <= 0.70128643;
cosLookup[8278] <= 0.701218076;
cosLookup[8279] <= 0.701149716;
cosLookup[8280] <= 0.701081349;
cosLookup[8281] <= 0.701012976;
cosLookup[8282] <= 0.700944596;
cosLookup[8283] <= 0.70087621;
cosLookup[8284] <= 0.700807818;
cosLookup[8285] <= 0.700739419;
cosLookup[8286] <= 0.700671013;
cosLookup[8287] <= 0.700602601;
cosLookup[8288] <= 0.700534183;
cosLookup[8289] <= 0.700465758;
cosLookup[8290] <= 0.700397327;
cosLookup[8291] <= 0.70032889;
cosLookup[8292] <= 0.700260445;
cosLookup[8293] <= 0.700191995;
cosLookup[8294] <= 0.700123538;
cosLookup[8295] <= 0.700055075;
cosLookup[8296] <= 0.699986605;
cosLookup[8297] <= 0.699918129;
cosLookup[8298] <= 0.699849646;
cosLookup[8299] <= 0.699781157;
cosLookup[8300] <= 0.699712661;
cosLookup[8301] <= 0.699644159;
cosLookup[8302] <= 0.699575651;
cosLookup[8303] <= 0.699507136;
cosLookup[8304] <= 0.699438615;
cosLookup[8305] <= 0.699370087;
cosLookup[8306] <= 0.699301553;
cosLookup[8307] <= 0.699233012;
cosLookup[8308] <= 0.699164465;
cosLookup[8309] <= 0.699095912;
cosLookup[8310] <= 0.699027352;
cosLookup[8311] <= 0.698958786;
cosLookup[8312] <= 0.698890213;
cosLookup[8313] <= 0.698821634;
cosLookup[8314] <= 0.698753049;
cosLookup[8315] <= 0.698684457;
cosLookup[8316] <= 0.698615858;
cosLookup[8317] <= 0.698547253;
cosLookup[8318] <= 0.698478642;
cosLookup[8319] <= 0.698410025;
cosLookup[8320] <= 0.6983414;
cosLookup[8321] <= 0.69827277;
cosLookup[8322] <= 0.698204133;
cosLookup[8323] <= 0.69813549;
cosLookup[8324] <= 0.69806684;
cosLookup[8325] <= 0.697998184;
cosLookup[8326] <= 0.697929521;
cosLookup[8327] <= 0.697860852;
cosLookup[8328] <= 0.697792177;
cosLookup[8329] <= 0.697723495;
cosLookup[8330] <= 0.697654807;
cosLookup[8331] <= 0.697586112;
cosLookup[8332] <= 0.697517411;
cosLookup[8333] <= 0.697448704;
cosLookup[8334] <= 0.69737999;
cosLookup[8335] <= 0.697311269;
cosLookup[8336] <= 0.697242543;
cosLookup[8337] <= 0.69717381;
cosLookup[8338] <= 0.69710507;
cosLookup[8339] <= 0.697036324;
cosLookup[8340] <= 0.696967572;
cosLookup[8341] <= 0.696898813;
cosLookup[8342] <= 0.696830048;
cosLookup[8343] <= 0.696761276;
cosLookup[8344] <= 0.696692498;
cosLookup[8345] <= 0.696623714;
cosLookup[8346] <= 0.696554923;
cosLookup[8347] <= 0.696486126;
cosLookup[8348] <= 0.696417322;
cosLookup[8349] <= 0.696348512;
cosLookup[8350] <= 0.696279696;
cosLookup[8351] <= 0.696210873;
cosLookup[8352] <= 0.696142044;
cosLookup[8353] <= 0.696073208;
cosLookup[8354] <= 0.696004366;
cosLookup[8355] <= 0.695935518;
cosLookup[8356] <= 0.695866663;
cosLookup[8357] <= 0.695797802;
cosLookup[8358] <= 0.695728934;
cosLookup[8359] <= 0.69566006;
cosLookup[8360] <= 0.69559118;
cosLookup[8361] <= 0.695522293;
cosLookup[8362] <= 0.6954534;
cosLookup[8363] <= 0.695384501;
cosLookup[8364] <= 0.695315595;
cosLookup[8365] <= 0.695246682;
cosLookup[8366] <= 0.695177764;
cosLookup[8367] <= 0.695108838;
cosLookup[8368] <= 0.695039907;
cosLookup[8369] <= 0.694970969;
cosLookup[8370] <= 0.694902025;
cosLookup[8371] <= 0.694833074;
cosLookup[8372] <= 0.694764117;
cosLookup[8373] <= 0.694695154;
cosLookup[8374] <= 0.694626184;
cosLookup[8375] <= 0.694557208;
cosLookup[8376] <= 0.694488225;
cosLookup[8377] <= 0.694419236;
cosLookup[8378] <= 0.694350241;
cosLookup[8379] <= 0.694281239;
cosLookup[8380] <= 0.694212231;
cosLookup[8381] <= 0.694143216;
cosLookup[8382] <= 0.694074195;
cosLookup[8383] <= 0.694005168;
cosLookup[8384] <= 0.693936134;
cosLookup[8385] <= 0.693867094;
cosLookup[8386] <= 0.693798048;
cosLookup[8387] <= 0.693728995;
cosLookup[8388] <= 0.693659936;
cosLookup[8389] <= 0.69359087;
cosLookup[8390] <= 0.693521798;
cosLookup[8391] <= 0.69345272;
cosLookup[8392] <= 0.693383635;
cosLookup[8393] <= 0.693314544;
cosLookup[8394] <= 0.693245447;
cosLookup[8395] <= 0.693176343;
cosLookup[8396] <= 0.693107233;
cosLookup[8397] <= 0.693038116;
cosLookup[8398] <= 0.692968993;
cosLookup[8399] <= 0.692899864;
cosLookup[8400] <= 0.692830728;
cosLookup[8401] <= 0.692761586;
cosLookup[8402] <= 0.692692438;
cosLookup[8403] <= 0.692623283;
cosLookup[8404] <= 0.692554122;
cosLookup[8405] <= 0.692484955;
cosLookup[8406] <= 0.692415781;
cosLookup[8407] <= 0.692346601;
cosLookup[8408] <= 0.692277414;
cosLookup[8409] <= 0.692208221;
cosLookup[8410] <= 0.692139022;
cosLookup[8411] <= 0.692069816;
cosLookup[8412] <= 0.692000604;
cosLookup[8413] <= 0.691931386;
cosLookup[8414] <= 0.691862161;
cosLookup[8415] <= 0.69179293;
cosLookup[8416] <= 0.691723692;
cosLookup[8417] <= 0.691654448;
cosLookup[8418] <= 0.691585198;
cosLookup[8419] <= 0.691515942;
cosLookup[8420] <= 0.691446679;
cosLookup[8421] <= 0.691377409;
cosLookup[8422] <= 0.691308134;
cosLookup[8423] <= 0.691238852;
cosLookup[8424] <= 0.691169563;
cosLookup[8425] <= 0.691100269;
cosLookup[8426] <= 0.691030968;
cosLookup[8427] <= 0.69096166;
cosLookup[8428] <= 0.690892347;
cosLookup[8429] <= 0.690823026;
cosLookup[8430] <= 0.6907537;
cosLookup[8431] <= 0.690684367;
cosLookup[8432] <= 0.690615028;
cosLookup[8433] <= 0.690545683;
cosLookup[8434] <= 0.690476331;
cosLookup[8435] <= 0.690406973;
cosLookup[8436] <= 0.690337608;
cosLookup[8437] <= 0.690268237;
cosLookup[8438] <= 0.69019886;
cosLookup[8439] <= 0.690129476;
cosLookup[8440] <= 0.690060086;
cosLookup[8441] <= 0.68999069;
cosLookup[8442] <= 0.689921287;
cosLookup[8443] <= 0.689851878;
cosLookup[8444] <= 0.689782463;
cosLookup[8445] <= 0.689713042;
cosLookup[8446] <= 0.689643614;
cosLookup[8447] <= 0.689574179;
cosLookup[8448] <= 0.689504739;
cosLookup[8449] <= 0.689435292;
cosLookup[8450] <= 0.689365838;
cosLookup[8451] <= 0.689296379;
cosLookup[8452] <= 0.689226913;
cosLookup[8453] <= 0.68915744;
cosLookup[8454] <= 0.689087962;
cosLookup[8455] <= 0.689018477;
cosLookup[8456] <= 0.688948985;
cosLookup[8457] <= 0.688879488;
cosLookup[8458] <= 0.688809984;
cosLookup[8459] <= 0.688740473;
cosLookup[8460] <= 0.688670957;
cosLookup[8461] <= 0.688601433;
cosLookup[8462] <= 0.688531904;
cosLookup[8463] <= 0.688462368;
cosLookup[8464] <= 0.688392826;
cosLookup[8465] <= 0.688323278;
cosLookup[8466] <= 0.688253724;
cosLookup[8467] <= 0.688184163;
cosLookup[8468] <= 0.688114595;
cosLookup[8469] <= 0.688045022;
cosLookup[8470] <= 0.687975442;
cosLookup[8471] <= 0.687905855;
cosLookup[8472] <= 0.687836263;
cosLookup[8473] <= 0.687766664;
cosLookup[8474] <= 0.687697059;
cosLookup[8475] <= 0.687627447;
cosLookup[8476] <= 0.687557829;
cosLookup[8477] <= 0.687488205;
cosLookup[8478] <= 0.687418574;
cosLookup[8479] <= 0.687348937;
cosLookup[8480] <= 0.687279294;
cosLookup[8481] <= 0.687209645;
cosLookup[8482] <= 0.687139989;
cosLookup[8483] <= 0.687070327;
cosLookup[8484] <= 0.687000658;
cosLookup[8485] <= 0.686930984;
cosLookup[8486] <= 0.686861303;
cosLookup[8487] <= 0.686791615;
cosLookup[8488] <= 0.686721922;
cosLookup[8489] <= 0.686652222;
cosLookup[8490] <= 0.686582515;
cosLookup[8491] <= 0.686512803;
cosLookup[8492] <= 0.686443084;
cosLookup[8493] <= 0.686373358;
cosLookup[8494] <= 0.686303627;
cosLookup[8495] <= 0.686233889;
cosLookup[8496] <= 0.686164145;
cosLookup[8497] <= 0.686094394;
cosLookup[8498] <= 0.686024637;
cosLookup[8499] <= 0.685954874;
cosLookup[8500] <= 0.685885105;
cosLookup[8501] <= 0.685815329;
cosLookup[8502] <= 0.685745547;
cosLookup[8503] <= 0.685675759;
cosLookup[8504] <= 0.685605964;
cosLookup[8505] <= 0.685536163;
cosLookup[8506] <= 0.685466356;
cosLookup[8507] <= 0.685396542;
cosLookup[8508] <= 0.685326723;
cosLookup[8509] <= 0.685256897;
cosLookup[8510] <= 0.685187064;
cosLookup[8511] <= 0.685117225;
cosLookup[8512] <= 0.68504738;
cosLookup[8513] <= 0.684977529;
cosLookup[8514] <= 0.684907671;
cosLookup[8515] <= 0.684837807;
cosLookup[8516] <= 0.684767937;
cosLookup[8517] <= 0.684698061;
cosLookup[8518] <= 0.684628178;
cosLookup[8519] <= 0.684558289;
cosLookup[8520] <= 0.684488393;
cosLookup[8521] <= 0.684418492;
cosLookup[8522] <= 0.684348584;
cosLookup[8523] <= 0.684278669;
cosLookup[8524] <= 0.684208749;
cosLookup[8525] <= 0.684138822;
cosLookup[8526] <= 0.684068889;
cosLookup[8527] <= 0.683998949;
cosLookup[8528] <= 0.683929004;
cosLookup[8529] <= 0.683859052;
cosLookup[8530] <= 0.683789093;
cosLookup[8531] <= 0.683719129;
cosLookup[8532] <= 0.683649158;
cosLookup[8533] <= 0.683579181;
cosLookup[8534] <= 0.683509197;
cosLookup[8535] <= 0.683439208;
cosLookup[8536] <= 0.683369212;
cosLookup[8537] <= 0.683299209;
cosLookup[8538] <= 0.683229201;
cosLookup[8539] <= 0.683159186;
cosLookup[8540] <= 0.683089165;
cosLookup[8541] <= 0.683019137;
cosLookup[8542] <= 0.682949104;
cosLookup[8543] <= 0.682879064;
cosLookup[8544] <= 0.682809018;
cosLookup[8545] <= 0.682738965;
cosLookup[8546] <= 0.682668906;
cosLookup[8547] <= 0.682598841;
cosLookup[8548] <= 0.68252877;
cosLookup[8549] <= 0.682458692;
cosLookup[8550] <= 0.682388608;
cosLookup[8551] <= 0.682318518;
cosLookup[8552] <= 0.682248422;
cosLookup[8553] <= 0.682178319;
cosLookup[8554] <= 0.68210821;
cosLookup[8555] <= 0.682038095;
cosLookup[8556] <= 0.681967973;
cosLookup[8557] <= 0.681897846;
cosLookup[8558] <= 0.681827711;
cosLookup[8559] <= 0.681757571;
cosLookup[8560] <= 0.681687425;
cosLookup[8561] <= 0.681617272;
cosLookup[8562] <= 0.681547113;
cosLookup[8563] <= 0.681476947;
cosLookup[8564] <= 0.681406776;
cosLookup[8565] <= 0.681336598;
cosLookup[8566] <= 0.681266413;
cosLookup[8567] <= 0.681196223;
cosLookup[8568] <= 0.681126026;
cosLookup[8569] <= 0.681055823;
cosLookup[8570] <= 0.680985614;
cosLookup[8571] <= 0.680915399;
cosLookup[8572] <= 0.680845177;
cosLookup[8573] <= 0.680774949;
cosLookup[8574] <= 0.680704715;
cosLookup[8575] <= 0.680634474;
cosLookup[8576] <= 0.680564227;
cosLookup[8577] <= 0.680493974;
cosLookup[8578] <= 0.680423715;
cosLookup[8579] <= 0.680353449;
cosLookup[8580] <= 0.680283178;
cosLookup[8581] <= 0.680212899;
cosLookup[8582] <= 0.680142615;
cosLookup[8583] <= 0.680072325;
cosLookup[8584] <= 0.680002028;
cosLookup[8585] <= 0.679931725;
cosLookup[8586] <= 0.679861415;
cosLookup[8587] <= 0.6797911;
cosLookup[8588] <= 0.679720778;
cosLookup[8589] <= 0.67965045;
cosLookup[8590] <= 0.679580116;
cosLookup[8591] <= 0.679509775;
cosLookup[8592] <= 0.679439428;
cosLookup[8593] <= 0.679369075;
cosLookup[8594] <= 0.679298716;
cosLookup[8595] <= 0.67922835;
cosLookup[8596] <= 0.679157979;
cosLookup[8597] <= 0.679087601;
cosLookup[8598] <= 0.679017216;
cosLookup[8599] <= 0.678946826;
cosLookup[8600] <= 0.678876429;
cosLookup[8601] <= 0.678806026;
cosLookup[8602] <= 0.678735617;
cosLookup[8603] <= 0.678665201;
cosLookup[8604] <= 0.67859478;
cosLookup[8605] <= 0.678524352;
cosLookup[8606] <= 0.678453917;
cosLookup[8607] <= 0.678383477;
cosLookup[8608] <= 0.67831303;
cosLookup[8609] <= 0.678242577;
cosLookup[8610] <= 0.678172118;
cosLookup[8611] <= 0.678101653;
cosLookup[8612] <= 0.678031181;
cosLookup[8613] <= 0.677960703;
cosLookup[8614] <= 0.677890219;
cosLookup[8615] <= 0.677819729;
cosLookup[8616] <= 0.677749233;
cosLookup[8617] <= 0.67767873;
cosLookup[8618] <= 0.677608221;
cosLookup[8619] <= 0.677537706;
cosLookup[8620] <= 0.677467184;
cosLookup[8621] <= 0.677396656;
cosLookup[8622] <= 0.677326123;
cosLookup[8623] <= 0.677255582;
cosLookup[8624] <= 0.677185036;
cosLookup[8625] <= 0.677114483;
cosLookup[8626] <= 0.677043925;
cosLookup[8627] <= 0.67697336;
cosLookup[8628] <= 0.676902788;
cosLookup[8629] <= 0.676832211;
cosLookup[8630] <= 0.676761627;
cosLookup[8631] <= 0.676691037;
cosLookup[8632] <= 0.676620441;
cosLookup[8633] <= 0.676549839;
cosLookup[8634] <= 0.67647923;
cosLookup[8635] <= 0.676408615;
cosLookup[8636] <= 0.676337994;
cosLookup[8637] <= 0.676267367;
cosLookup[8638] <= 0.676196734;
cosLookup[8639] <= 0.676126094;
cosLookup[8640] <= 0.676055448;
cosLookup[8641] <= 0.675984796;
cosLookup[8642] <= 0.675914138;
cosLookup[8643] <= 0.675843473;
cosLookup[8644] <= 0.675772802;
cosLookup[8645] <= 0.675702125;
cosLookup[8646] <= 0.675631442;
cosLookup[8647] <= 0.675560753;
cosLookup[8648] <= 0.675490057;
cosLookup[8649] <= 0.675419356;
cosLookup[8650] <= 0.675348648;
cosLookup[8651] <= 0.675277933;
cosLookup[8652] <= 0.675207213;
cosLookup[8653] <= 0.675136486;
cosLookup[8654] <= 0.675065753;
cosLookup[8655] <= 0.674995014;
cosLookup[8656] <= 0.674924269;
cosLookup[8657] <= 0.674853518;
cosLookup[8658] <= 0.67478276;
cosLookup[8659] <= 0.674711996;
cosLookup[8660] <= 0.674641226;
cosLookup[8661] <= 0.67457045;
cosLookup[8662] <= 0.674499667;
cosLookup[8663] <= 0.674428879;
cosLookup[8664] <= 0.674358084;
cosLookup[8665] <= 0.674287283;
cosLookup[8666] <= 0.674216476;
cosLookup[8667] <= 0.674145662;
cosLookup[8668] <= 0.674074842;
cosLookup[8669] <= 0.674004017;
cosLookup[8670] <= 0.673933185;
cosLookup[8671] <= 0.673862346;
cosLookup[8672] <= 0.673791502;
cosLookup[8673] <= 0.673720651;
cosLookup[8674] <= 0.673649794;
cosLookup[8675] <= 0.673578931;
cosLookup[8676] <= 0.673508062;
cosLookup[8677] <= 0.673437187;
cosLookup[8678] <= 0.673366305;
cosLookup[8679] <= 0.673295417;
cosLookup[8680] <= 0.673224523;
cosLookup[8681] <= 0.673153623;
cosLookup[8682] <= 0.673082717;
cosLookup[8683] <= 0.673011804;
cosLookup[8684] <= 0.672940886;
cosLookup[8685] <= 0.672869961;
cosLookup[8686] <= 0.67279903;
cosLookup[8687] <= 0.672728092;
cosLookup[8688] <= 0.672657149;
cosLookup[8689] <= 0.672586199;
cosLookup[8690] <= 0.672515243;
cosLookup[8691] <= 0.672444281;
cosLookup[8692] <= 0.672373313;
cosLookup[8693] <= 0.672302339;
cosLookup[8694] <= 0.672231358;
cosLookup[8695] <= 0.672160371;
cosLookup[8696] <= 0.672089379;
cosLookup[8697] <= 0.672018379;
cosLookup[8698] <= 0.671947374;
cosLookup[8699] <= 0.671876363;
cosLookup[8700] <= 0.671805345;
cosLookup[8701] <= 0.671734321;
cosLookup[8702] <= 0.671663291;
cosLookup[8703] <= 0.671592255;
cosLookup[8704] <= 0.671521213;
cosLookup[8705] <= 0.671450164;
cosLookup[8706] <= 0.67137911;
cosLookup[8707] <= 0.671308049;
cosLookup[8708] <= 0.671236982;
cosLookup[8709] <= 0.671165909;
cosLookup[8710] <= 0.671094829;
cosLookup[8711] <= 0.671023744;
cosLookup[8712] <= 0.670952652;
cosLookup[8713] <= 0.670881554;
cosLookup[8714] <= 0.67081045;
cosLookup[8715] <= 0.67073934;
cosLookup[8716] <= 0.670668224;
cosLookup[8717] <= 0.670597101;
cosLookup[8718] <= 0.670525972;
cosLookup[8719] <= 0.670454837;
cosLookup[8720] <= 0.670383696;
cosLookup[8721] <= 0.670312549;
cosLookup[8722] <= 0.670241396;
cosLookup[8723] <= 0.670170236;
cosLookup[8724] <= 0.670099071;
cosLookup[8725] <= 0.670027899;
cosLookup[8726] <= 0.669956721;
cosLookup[8727] <= 0.669885537;
cosLookup[8728] <= 0.669814346;
cosLookup[8729] <= 0.66974315;
cosLookup[8730] <= 0.669671947;
cosLookup[8731] <= 0.669600739;
cosLookup[8732] <= 0.669529524;
cosLookup[8733] <= 0.669458303;
cosLookup[8734] <= 0.669387075;
cosLookup[8735] <= 0.669315842;
cosLookup[8736] <= 0.669244602;
cosLookup[8737] <= 0.669173357;
cosLookup[8738] <= 0.669102105;
cosLookup[8739] <= 0.669030847;
cosLookup[8740] <= 0.668959583;
cosLookup[8741] <= 0.668888312;
cosLookup[8742] <= 0.668817036;
cosLookup[8743] <= 0.668745753;
cosLookup[8744] <= 0.668674465;
cosLookup[8745] <= 0.66860317;
cosLookup[8746] <= 0.668531869;
cosLookup[8747] <= 0.668460561;
cosLookup[8748] <= 0.668389248;
cosLookup[8749] <= 0.668317929;
cosLookup[8750] <= 0.668246603;
cosLookup[8751] <= 0.668175271;
cosLookup[8752] <= 0.668103933;
cosLookup[8753] <= 0.668032589;
cosLookup[8754] <= 0.667961239;
cosLookup[8755] <= 0.667889883;
cosLookup[8756] <= 0.66781852;
cosLookup[8757] <= 0.667747152;
cosLookup[8758] <= 0.667675777;
cosLookup[8759] <= 0.667604396;
cosLookup[8760] <= 0.667533009;
cosLookup[8761] <= 0.667461616;
cosLookup[8762] <= 0.667390217;
cosLookup[8763] <= 0.667318811;
cosLookup[8764] <= 0.6672474;
cosLookup[8765] <= 0.667175982;
cosLookup[8766] <= 0.667104558;
cosLookup[8767] <= 0.667033128;
cosLookup[8768] <= 0.666961692;
cosLookup[8769] <= 0.66689025;
cosLookup[8770] <= 0.666818801;
cosLookup[8771] <= 0.666747347;
cosLookup[8772] <= 0.666675886;
cosLookup[8773] <= 0.66660442;
cosLookup[8774] <= 0.666532947;
cosLookup[8775] <= 0.666461468;
cosLookup[8776] <= 0.666389983;
cosLookup[8777] <= 0.666318491;
cosLookup[8778] <= 0.666246994;
cosLookup[8779] <= 0.66617549;
cosLookup[8780] <= 0.666103981;
cosLookup[8781] <= 0.666032465;
cosLookup[8782] <= 0.665960943;
cosLookup[8783] <= 0.665889415;
cosLookup[8784] <= 0.665817881;
cosLookup[8785] <= 0.665746341;
cosLookup[8786] <= 0.665674795;
cosLookup[8787] <= 0.665603242;
cosLookup[8788] <= 0.665531683;
cosLookup[8789] <= 0.665460119;
cosLookup[8790] <= 0.665388548;
cosLookup[8791] <= 0.665316971;
cosLookup[8792] <= 0.665245388;
cosLookup[8793] <= 0.665173799;
cosLookup[8794] <= 0.665102203;
cosLookup[8795] <= 0.665030602;
cosLookup[8796] <= 0.664958994;
cosLookup[8797] <= 0.664887381;
cosLookup[8798] <= 0.664815761;
cosLookup[8799] <= 0.664744135;
cosLookup[8800] <= 0.664672503;
cosLookup[8801] <= 0.664600865;
cosLookup[8802] <= 0.664529221;
cosLookup[8803] <= 0.664457571;
cosLookup[8804] <= 0.664385914;
cosLookup[8805] <= 0.664314252;
cosLookup[8806] <= 0.664242583;
cosLookup[8807] <= 0.664170908;
cosLookup[8808] <= 0.664099228;
cosLookup[8809] <= 0.664027541;
cosLookup[8810] <= 0.663955848;
cosLookup[8811] <= 0.663884148;
cosLookup[8812] <= 0.663812443;
cosLookup[8813] <= 0.663740732;
cosLookup[8814] <= 0.663669014;
cosLookup[8815] <= 0.663597291;
cosLookup[8816] <= 0.663525561;
cosLookup[8817] <= 0.663453825;
cosLookup[8818] <= 0.663382084;
cosLookup[8819] <= 0.663310336;
cosLookup[8820] <= 0.663238582;
cosLookup[8821] <= 0.663166821;
cosLookup[8822] <= 0.663095055;
cosLookup[8823] <= 0.663023283;
cosLookup[8824] <= 0.662951504;
cosLookup[8825] <= 0.66287972;
cosLookup[8826] <= 0.662807929;
cosLookup[8827] <= 0.662736132;
cosLookup[8828] <= 0.66266433;
cosLookup[8829] <= 0.662592521;
cosLookup[8830] <= 0.662520706;
cosLookup[8831] <= 0.662448885;
cosLookup[8832] <= 0.662377057;
cosLookup[8833] <= 0.662305224;
cosLookup[8834] <= 0.662233385;
cosLookup[8835] <= 0.662161539;
cosLookup[8836] <= 0.662089688;
cosLookup[8837] <= 0.66201783;
cosLookup[8838] <= 0.661945967;
cosLookup[8839] <= 0.661874097;
cosLookup[8840] <= 0.661802221;
cosLookup[8841] <= 0.661730339;
cosLookup[8842] <= 0.661658451;
cosLookup[8843] <= 0.661586557;
cosLookup[8844] <= 0.661514657;
cosLookup[8845] <= 0.66144275;
cosLookup[8846] <= 0.661370838;
cosLookup[8847] <= 0.66129892;
cosLookup[8848] <= 0.661226995;
cosLookup[8849] <= 0.661155064;
cosLookup[8850] <= 0.661083128;
cosLookup[8851] <= 0.661011185;
cosLookup[8852] <= 0.660939236;
cosLookup[8853] <= 0.660867281;
cosLookup[8854] <= 0.66079532;
cosLookup[8855] <= 0.660723353;
cosLookup[8856] <= 0.66065138;
cosLookup[8857] <= 0.660579401;
cosLookup[8858] <= 0.660507416;
cosLookup[8859] <= 0.660435424;
cosLookup[8860] <= 0.660363427;
cosLookup[8861] <= 0.660291423;
cosLookup[8862] <= 0.660219414;
cosLookup[8863] <= 0.660147398;
cosLookup[8864] <= 0.660075376;
cosLookup[8865] <= 0.660003349;
cosLookup[8866] <= 0.659931315;
cosLookup[8867] <= 0.659859275;
cosLookup[8868] <= 0.659787229;
cosLookup[8869] <= 0.659715177;
cosLookup[8870] <= 0.659643119;
cosLookup[8871] <= 0.659571055;
cosLookup[8872] <= 0.659498984;
cosLookup[8873] <= 0.659426908;
cosLookup[8874] <= 0.659354826;
cosLookup[8875] <= 0.659282737;
cosLookup[8876] <= 0.659210643;
cosLookup[8877] <= 0.659138542;
cosLookup[8878] <= 0.659066436;
cosLookup[8879] <= 0.658994323;
cosLookup[8880] <= 0.658922204;
cosLookup[8881] <= 0.65885008;
cosLookup[8882] <= 0.658777949;
cosLookup[8883] <= 0.658705812;
cosLookup[8884] <= 0.658633669;
cosLookup[8885] <= 0.65856152;
cosLookup[8886] <= 0.658489365;
cosLookup[8887] <= 0.658417204;
cosLookup[8888] <= 0.658345037;
cosLookup[8889] <= 0.658272864;
cosLookup[8890] <= 0.658200684;
cosLookup[8891] <= 0.658128499;
cosLookup[8892] <= 0.658056308;
cosLookup[8893] <= 0.65798411;
cosLookup[8894] <= 0.657911907;
cosLookup[8895] <= 0.657839697;
cosLookup[8896] <= 0.657767482;
cosLookup[8897] <= 0.65769526;
cosLookup[8898] <= 0.657623033;
cosLookup[8899] <= 0.657550799;
cosLookup[8900] <= 0.657478559;
cosLookup[8901] <= 0.657406313;
cosLookup[8902] <= 0.657334062;
cosLookup[8903] <= 0.657261804;
cosLookup[8904] <= 0.65718954;
cosLookup[8905] <= 0.65711727;
cosLookup[8906] <= 0.657044994;
cosLookup[8907] <= 0.656972712;
cosLookup[8908] <= 0.656900424;
cosLookup[8909] <= 0.65682813;
cosLookup[8910] <= 0.656755829;
cosLookup[8911] <= 0.656683523;
cosLookup[8912] <= 0.656611211;
cosLookup[8913] <= 0.656538893;
cosLookup[8914] <= 0.656466569;
cosLookup[8915] <= 0.656394238;
cosLookup[8916] <= 0.656321902;
cosLookup[8917] <= 0.656249559;
cosLookup[8918] <= 0.656177211;
cosLookup[8919] <= 0.656104857;
cosLookup[8920] <= 0.656032496;
cosLookup[8921] <= 0.65596013;
cosLookup[8922] <= 0.655887757;
cosLookup[8923] <= 0.655815378;
cosLookup[8924] <= 0.655742994;
cosLookup[8925] <= 0.655670603;
cosLookup[8926] <= 0.655598207;
cosLookup[8927] <= 0.655525804;
cosLookup[8928] <= 0.655453395;
cosLookup[8929] <= 0.65538098;
cosLookup[8930] <= 0.65530856;
cosLookup[8931] <= 0.655236133;
cosLookup[8932] <= 0.6551637;
cosLookup[8933] <= 0.655091261;
cosLookup[8934] <= 0.655018816;
cosLookup[8935] <= 0.654946365;
cosLookup[8936] <= 0.654873909;
cosLookup[8937] <= 0.654801446;
cosLookup[8938] <= 0.654728977;
cosLookup[8939] <= 0.654656502;
cosLookup[8940] <= 0.654584021;
cosLookup[8941] <= 0.654511534;
cosLookup[8942] <= 0.654439041;
cosLookup[8943] <= 0.654366542;
cosLookup[8944] <= 0.654294037;
cosLookup[8945] <= 0.654221526;
cosLookup[8946] <= 0.654149009;
cosLookup[8947] <= 0.654076485;
cosLookup[8948] <= 0.654003956;
cosLookup[8949] <= 0.653931421;
cosLookup[8950] <= 0.65385888;
cosLookup[8951] <= 0.653786333;
cosLookup[8952] <= 0.65371378;
cosLookup[8953] <= 0.653641221;
cosLookup[8954] <= 0.653568656;
cosLookup[8955] <= 0.653496084;
cosLookup[8956] <= 0.653423507;
cosLookup[8957] <= 0.653350924;
cosLookup[8958] <= 0.653278335;
cosLookup[8959] <= 0.65320574;
cosLookup[8960] <= 0.653133138;
cosLookup[8961] <= 0.653060531;
cosLookup[8962] <= 0.652987918;
cosLookup[8963] <= 0.652915299;
cosLookup[8964] <= 0.652842674;
cosLookup[8965] <= 0.652770042;
cosLookup[8966] <= 0.652697405;
cosLookup[8967] <= 0.652624762;
cosLookup[8968] <= 0.652552113;
cosLookup[8969] <= 0.652479458;
cosLookup[8970] <= 0.652406796;
cosLookup[8971] <= 0.652334129;
cosLookup[8972] <= 0.652261456;
cosLookup[8973] <= 0.652188777;
cosLookup[8974] <= 0.652116091;
cosLookup[8975] <= 0.6520434;
cosLookup[8976] <= 0.651970703;
cosLookup[8977] <= 0.651898;
cosLookup[8978] <= 0.651825291;
cosLookup[8979] <= 0.651752576;
cosLookup[8980] <= 0.651679854;
cosLookup[8981] <= 0.651607127;
cosLookup[8982] <= 0.651534394;
cosLookup[8983] <= 0.651461655;
cosLookup[8984] <= 0.65138891;
cosLookup[8985] <= 0.651316159;
cosLookup[8986] <= 0.651243402;
cosLookup[8987] <= 0.651170639;
cosLookup[8988] <= 0.65109787;
cosLookup[8989] <= 0.651025094;
cosLookup[8990] <= 0.650952313;
cosLookup[8991] <= 0.650879526;
cosLookup[8992] <= 0.650806733;
cosLookup[8993] <= 0.650733934;
cosLookup[8994] <= 0.650661129;
cosLookup[8995] <= 0.650588319;
cosLookup[8996] <= 0.650515502;
cosLookup[8997] <= 0.650442679;
cosLookup[8998] <= 0.65036985;
cosLookup[8999] <= 0.650297015;
cosLookup[9000] <= 0.650224174;
cosLookup[9001] <= 0.650151327;
cosLookup[9002] <= 0.650078474;
cosLookup[9003] <= 0.650005616;
cosLookup[9004] <= 0.649932751;
cosLookup[9005] <= 0.64985988;
cosLookup[9006] <= 0.649787003;
cosLookup[9007] <= 0.649714121;
cosLookup[9008] <= 0.649641232;
cosLookup[9009] <= 0.649568338;
cosLookup[9010] <= 0.649495437;
cosLookup[9011] <= 0.64942253;
cosLookup[9012] <= 0.649349618;
cosLookup[9013] <= 0.649276699;
cosLookup[9014] <= 0.649203775;
cosLookup[9015] <= 0.649130844;
cosLookup[9016] <= 0.649057908;
cosLookup[9017] <= 0.648984966;
cosLookup[9018] <= 0.648912017;
cosLookup[9019] <= 0.648839063;
cosLookup[9020] <= 0.648766103;
cosLookup[9021] <= 0.648693136;
cosLookup[9022] <= 0.648620164;
cosLookup[9023] <= 0.648547186;
cosLookup[9024] <= 0.648474202;
cosLookup[9025] <= 0.648401212;
cosLookup[9026] <= 0.648328216;
cosLookup[9027] <= 0.648255214;
cosLookup[9028] <= 0.648182206;
cosLookup[9029] <= 0.648109192;
cosLookup[9030] <= 0.648036172;
cosLookup[9031] <= 0.647963146;
cosLookup[9032] <= 0.647890114;
cosLookup[9033] <= 0.647817077;
cosLookup[9034] <= 0.647744033;
cosLookup[9035] <= 0.647670983;
cosLookup[9036] <= 0.647597928;
cosLookup[9037] <= 0.647524866;
cosLookup[9038] <= 0.647451799;
cosLookup[9039] <= 0.647378725;
cosLookup[9040] <= 0.647305646;
cosLookup[9041] <= 0.64723256;
cosLookup[9042] <= 0.647159469;
cosLookup[9043] <= 0.647086372;
cosLookup[9044] <= 0.647013269;
cosLookup[9045] <= 0.646940159;
cosLookup[9046] <= 0.646867044;
cosLookup[9047] <= 0.646793923;
cosLookup[9048] <= 0.646720796;
cosLookup[9049] <= 0.646647663;
cosLookup[9050] <= 0.646574524;
cosLookup[9051] <= 0.64650138;
cosLookup[9052] <= 0.646428229;
cosLookup[9053] <= 0.646355072;
cosLookup[9054] <= 0.646281909;
cosLookup[9055] <= 0.646208741;
cosLookup[9056] <= 0.646135566;
cosLookup[9057] <= 0.646062386;
cosLookup[9058] <= 0.645989199;
cosLookup[9059] <= 0.645916007;
cosLookup[9060] <= 0.645842809;
cosLookup[9061] <= 0.645769604;
cosLookup[9062] <= 0.645696394;
cosLookup[9063] <= 0.645623178;
cosLookup[9064] <= 0.645549956;
cosLookup[9065] <= 0.645476728;
cosLookup[9066] <= 0.645403494;
cosLookup[9067] <= 0.645330254;
cosLookup[9068] <= 0.645257008;
cosLookup[9069] <= 0.645183757;
cosLookup[9070] <= 0.645110499;
cosLookup[9071] <= 0.645037235;
cosLookup[9072] <= 0.644963966;
cosLookup[9073] <= 0.644890691;
cosLookup[9074] <= 0.644817409;
cosLookup[9075] <= 0.644744122;
cosLookup[9076] <= 0.644670829;
cosLookup[9077] <= 0.644597529;
cosLookup[9078] <= 0.644524224;
cosLookup[9079] <= 0.644450913;
cosLookup[9080] <= 0.644377596;
cosLookup[9081] <= 0.644304274;
cosLookup[9082] <= 0.644230945;
cosLookup[9083] <= 0.64415761;
cosLookup[9084] <= 0.64408427;
cosLookup[9085] <= 0.644010923;
cosLookup[9086] <= 0.643937571;
cosLookup[9087] <= 0.643864212;
cosLookup[9088] <= 0.643790848;
cosLookup[9089] <= 0.643717478;
cosLookup[9090] <= 0.643644102;
cosLookup[9091] <= 0.64357072;
cosLookup[9092] <= 0.643497332;
cosLookup[9093] <= 0.643423938;
cosLookup[9094] <= 0.643350538;
cosLookup[9095] <= 0.643277132;
cosLookup[9096] <= 0.643203721;
cosLookup[9097] <= 0.643130303;
cosLookup[9098] <= 0.64305688;
cosLookup[9099] <= 0.64298345;
cosLookup[9100] <= 0.642910015;
cosLookup[9101] <= 0.642836574;
cosLookup[9102] <= 0.642763127;
cosLookup[9103] <= 0.642689674;
cosLookup[9104] <= 0.642616215;
cosLookup[9105] <= 0.64254275;
cosLookup[9106] <= 0.642469279;
cosLookup[9107] <= 0.642395803;
cosLookup[9108] <= 0.64232232;
cosLookup[9109] <= 0.642248832;
cosLookup[9110] <= 0.642175337;
cosLookup[9111] <= 0.642101837;
cosLookup[9112] <= 0.642028331;
cosLookup[9113] <= 0.641954819;
cosLookup[9114] <= 0.641881301;
cosLookup[9115] <= 0.641807777;
cosLookup[9116] <= 0.641734247;
cosLookup[9117] <= 0.641660712;
cosLookup[9118] <= 0.64158717;
cosLookup[9119] <= 0.641513623;
cosLookup[9120] <= 0.641440069;
cosLookup[9121] <= 0.64136651;
cosLookup[9122] <= 0.641292945;
cosLookup[9123] <= 0.641219374;
cosLookup[9124] <= 0.641145797;
cosLookup[9125] <= 0.641072214;
cosLookup[9126] <= 0.640998625;
cosLookup[9127] <= 0.640925031;
cosLookup[9128] <= 0.64085143;
cosLookup[9129] <= 0.640777824;
cosLookup[9130] <= 0.640704212;
cosLookup[9131] <= 0.640630593;
cosLookup[9132] <= 0.640556969;
cosLookup[9133] <= 0.640483339;
cosLookup[9134] <= 0.640409704;
cosLookup[9135] <= 0.640336062;
cosLookup[9136] <= 0.640262414;
cosLookup[9137] <= 0.640188761;
cosLookup[9138] <= 0.640115101;
cosLookup[9139] <= 0.640041436;
cosLookup[9140] <= 0.639967765;
cosLookup[9141] <= 0.639894088;
cosLookup[9142] <= 0.639820405;
cosLookup[9143] <= 0.639746716;
cosLookup[9144] <= 0.639673022;
cosLookup[9145] <= 0.639599321;
cosLookup[9146] <= 0.639525615;
cosLookup[9147] <= 0.639451902;
cosLookup[9148] <= 0.639378184;
cosLookup[9149] <= 0.63930446;
cosLookup[9150] <= 0.63923073;
cosLookup[9151] <= 0.639156994;
cosLookup[9152] <= 0.639083252;
cosLookup[9153] <= 0.639009505;
cosLookup[9154] <= 0.638935751;
cosLookup[9155] <= 0.638861992;
cosLookup[9156] <= 0.638788227;
cosLookup[9157] <= 0.638714456;
cosLookup[9158] <= 0.638640679;
cosLookup[9159] <= 0.638566896;
cosLookup[9160] <= 0.638493107;
cosLookup[9161] <= 0.638419313;
cosLookup[9162] <= 0.638345512;
cosLookup[9163] <= 0.638271706;
cosLookup[9164] <= 0.638197894;
cosLookup[9165] <= 0.638124076;
cosLookup[9166] <= 0.638050252;
cosLookup[9167] <= 0.637976422;
cosLookup[9168] <= 0.637902587;
cosLookup[9169] <= 0.637828745;
cosLookup[9170] <= 0.637754898;
cosLookup[9171] <= 0.637681045;
cosLookup[9172] <= 0.637607186;
cosLookup[9173] <= 0.637533321;
cosLookup[9174] <= 0.63745945;
cosLookup[9175] <= 0.637385573;
cosLookup[9176] <= 0.637311691;
cosLookup[9177] <= 0.637237802;
cosLookup[9178] <= 0.637163908;
cosLookup[9179] <= 0.637090008;
cosLookup[9180] <= 0.637016102;
cosLookup[9181] <= 0.63694219;
cosLookup[9182] <= 0.636868273;
cosLookup[9183] <= 0.636794349;
cosLookup[9184] <= 0.63672042;
cosLookup[9185] <= 0.636646484;
cosLookup[9186] <= 0.636572543;
cosLookup[9187] <= 0.636498596;
cosLookup[9188] <= 0.636424644;
cosLookup[9189] <= 0.636350685;
cosLookup[9190] <= 0.636276721;
cosLookup[9191] <= 0.63620275;
cosLookup[9192] <= 0.636128774;
cosLookup[9193] <= 0.636054792;
cosLookup[9194] <= 0.635980804;
cosLookup[9195] <= 0.63590681;
cosLookup[9196] <= 0.635832811;
cosLookup[9197] <= 0.635758805;
cosLookup[9198] <= 0.635684794;
cosLookup[9199] <= 0.635610777;
cosLookup[9200] <= 0.635536754;
cosLookup[9201] <= 0.635462725;
cosLookup[9202] <= 0.635388691;
cosLookup[9203] <= 0.63531465;
cosLookup[9204] <= 0.635240604;
cosLookup[9205] <= 0.635166552;
cosLookup[9206] <= 0.635092494;
cosLookup[9207] <= 0.63501843;
cosLookup[9208] <= 0.63494436;
cosLookup[9209] <= 0.634870285;
cosLookup[9210] <= 0.634796204;
cosLookup[9211] <= 0.634722116;
cosLookup[9212] <= 0.634648023;
cosLookup[9213] <= 0.634573925;
cosLookup[9214] <= 0.63449982;
cosLookup[9215] <= 0.634425709;
cosLookup[9216] <= 0.634351593;
cosLookup[9217] <= 0.634277471;
cosLookup[9218] <= 0.634203343;
cosLookup[9219] <= 0.634129209;
cosLookup[9220] <= 0.634055069;
cosLookup[9221] <= 0.633980924;
cosLookup[9222] <= 0.633906773;
cosLookup[9223] <= 0.633832615;
cosLookup[9224] <= 0.633758452;
cosLookup[9225] <= 0.633684284;
cosLookup[9226] <= 0.633610109;
cosLookup[9227] <= 0.633535929;
cosLookup[9228] <= 0.633461742;
cosLookup[9229] <= 0.63338755;
cosLookup[9230] <= 0.633313352;
cosLookup[9231] <= 0.633239149;
cosLookup[9232] <= 0.633164939;
cosLookup[9233] <= 0.633090724;
cosLookup[9234] <= 0.633016502;
cosLookup[9235] <= 0.632942275;
cosLookup[9236] <= 0.632868043;
cosLookup[9237] <= 0.632793804;
cosLookup[9238] <= 0.632719559;
cosLookup[9239] <= 0.632645309;
cosLookup[9240] <= 0.632571053;
cosLookup[9241] <= 0.632496791;
cosLookup[9242] <= 0.632422523;
cosLookup[9243] <= 0.63234825;
cosLookup[9244] <= 0.63227397;
cosLookup[9245] <= 0.632199685;
cosLookup[9246] <= 0.632125394;
cosLookup[9247] <= 0.632051097;
cosLookup[9248] <= 0.631976795;
cosLookup[9249] <= 0.631902486;
cosLookup[9250] <= 0.631828172;
cosLookup[9251] <= 0.631753852;
cosLookup[9252] <= 0.631679526;
cosLookup[9253] <= 0.631605195;
cosLookup[9254] <= 0.631530857;
cosLookup[9255] <= 0.631456514;
cosLookup[9256] <= 0.631382165;
cosLookup[9257] <= 0.63130781;
cosLookup[9258] <= 0.631233449;
cosLookup[9259] <= 0.631159083;
cosLookup[9260] <= 0.631084711;
cosLookup[9261] <= 0.631010333;
cosLookup[9262] <= 0.630935949;
cosLookup[9263] <= 0.630861559;
cosLookup[9264] <= 0.630787164;
cosLookup[9265] <= 0.630712762;
cosLookup[9266] <= 0.630638355;
cosLookup[9267] <= 0.630563942;
cosLookup[9268] <= 0.630489524;
cosLookup[9269] <= 0.630415099;
cosLookup[9270] <= 0.630340669;
cosLookup[9271] <= 0.630266233;
cosLookup[9272] <= 0.630191791;
cosLookup[9273] <= 0.630117343;
cosLookup[9274] <= 0.63004289;
cosLookup[9275] <= 0.629968431;
cosLookup[9276] <= 0.629893966;
cosLookup[9277] <= 0.629819495;
cosLookup[9278] <= 0.629745018;
cosLookup[9279] <= 0.629670536;
cosLookup[9280] <= 0.629596048;
cosLookup[9281] <= 0.629521554;
cosLookup[9282] <= 0.629447054;
cosLookup[9283] <= 0.629372548;
cosLookup[9284] <= 0.629298037;
cosLookup[9285] <= 0.62922352;
cosLookup[9286] <= 0.629148997;
cosLookup[9287] <= 0.629074468;
cosLookup[9288] <= 0.628999934;
cosLookup[9289] <= 0.628925394;
cosLookup[9290] <= 0.628850848;
cosLookup[9291] <= 0.628776296;
cosLookup[9292] <= 0.628701738;
cosLookup[9293] <= 0.628627175;
cosLookup[9294] <= 0.628552606;
cosLookup[9295] <= 0.628478031;
cosLookup[9296] <= 0.62840345;
cosLookup[9297] <= 0.628328864;
cosLookup[9298] <= 0.628254271;
cosLookup[9299] <= 0.628179673;
cosLookup[9300] <= 0.62810507;
cosLookup[9301] <= 0.62803046;
cosLookup[9302] <= 0.627955845;
cosLookup[9303] <= 0.627881223;
cosLookup[9304] <= 0.627806597;
cosLookup[9305] <= 0.627731964;
cosLookup[9306] <= 0.627657325;
cosLookup[9307] <= 0.627582681;
cosLookup[9308] <= 0.627508031;
cosLookup[9309] <= 0.627433376;
cosLookup[9310] <= 0.627358714;
cosLookup[9311] <= 0.627284047;
cosLookup[9312] <= 0.627209374;
cosLookup[9313] <= 0.627134695;
cosLookup[9314] <= 0.62706001;
cosLookup[9315] <= 0.62698532;
cosLookup[9316] <= 0.626910624;
cosLookup[9317] <= 0.626835922;
cosLookup[9318] <= 0.626761214;
cosLookup[9319] <= 0.626686501;
cosLookup[9320] <= 0.626611782;
cosLookup[9321] <= 0.626537057;
cosLookup[9322] <= 0.626462326;
cosLookup[9323] <= 0.62638759;
cosLookup[9324] <= 0.626312848;
cosLookup[9325] <= 0.6262381;
cosLookup[9326] <= 0.626163346;
cosLookup[9327] <= 0.626088586;
cosLookup[9328] <= 0.626013821;
cosLookup[9329] <= 0.62593905;
cosLookup[9330] <= 0.625864273;
cosLookup[9331] <= 0.625789491;
cosLookup[9332] <= 0.625714703;
cosLookup[9333] <= 0.625639909;
cosLookup[9334] <= 0.625565109;
cosLookup[9335] <= 0.625490304;
cosLookup[9336] <= 0.625415492;
cosLookup[9337] <= 0.625340675;
cosLookup[9338] <= 0.625265853;
cosLookup[9339] <= 0.625191024;
cosLookup[9340] <= 0.62511619;
cosLookup[9341] <= 0.62504135;
cosLookup[9342] <= 0.624966504;
cosLookup[9343] <= 0.624891653;
cosLookup[9344] <= 0.624816795;
cosLookup[9345] <= 0.624741932;
cosLookup[9346] <= 0.624667064;
cosLookup[9347] <= 0.624592189;
cosLookup[9348] <= 0.624517309;
cosLookup[9349] <= 0.624442423;
cosLookup[9350] <= 0.624367532;
cosLookup[9351] <= 0.624292634;
cosLookup[9352] <= 0.624217731;
cosLookup[9353] <= 0.624142822;
cosLookup[9354] <= 0.624067907;
cosLookup[9355] <= 0.623992987;
cosLookup[9356] <= 0.623918061;
cosLookup[9357] <= 0.623843129;
cosLookup[9358] <= 0.623768192;
cosLookup[9359] <= 0.623693248;
cosLookup[9360] <= 0.623618299;
cosLookup[9361] <= 0.623543344;
cosLookup[9362] <= 0.623468384;
cosLookup[9363] <= 0.623393418;
cosLookup[9364] <= 0.623318446;
cosLookup[9365] <= 0.623243468;
cosLookup[9366] <= 0.623168485;
cosLookup[9367] <= 0.623093496;
cosLookup[9368] <= 0.623018501;
cosLookup[9369] <= 0.6229435;
cosLookup[9370] <= 0.622868494;
cosLookup[9371] <= 0.622793482;
cosLookup[9372] <= 0.622718464;
cosLookup[9373] <= 0.62264344;
cosLookup[9374] <= 0.622568411;
cosLookup[9375] <= 0.622493376;
cosLookup[9376] <= 0.622418335;
cosLookup[9377] <= 0.622343289;
cosLookup[9378] <= 0.622268237;
cosLookup[9379] <= 0.622193179;
cosLookup[9380] <= 0.622118116;
cosLookup[9381] <= 0.622043046;
cosLookup[9382] <= 0.621967971;
cosLookup[9383] <= 0.621892891;
cosLookup[9384] <= 0.621817804;
cosLookup[9385] <= 0.621742712;
cosLookup[9386] <= 0.621667614;
cosLookup[9387] <= 0.621592511;
cosLookup[9388] <= 0.621517401;
cosLookup[9389] <= 0.621442286;
cosLookup[9390] <= 0.621367165;
cosLookup[9391] <= 0.621292039;
cosLookup[9392] <= 0.621216907;
cosLookup[9393] <= 0.621141769;
cosLookup[9394] <= 0.621066625;
cosLookup[9395] <= 0.620991476;
cosLookup[9396] <= 0.620916321;
cosLookup[9397] <= 0.620841161;
cosLookup[9398] <= 0.620765994;
cosLookup[9399] <= 0.620690822;
cosLookup[9400] <= 0.620615644;
cosLookup[9401] <= 0.620540461;
cosLookup[9402] <= 0.620465271;
cosLookup[9403] <= 0.620390077;
cosLookup[9404] <= 0.620314876;
cosLookup[9405] <= 0.62023967;
cosLookup[9406] <= 0.620164458;
cosLookup[9407] <= 0.62008924;
cosLookup[9408] <= 0.620014016;
cosLookup[9409] <= 0.619938787;
cosLookup[9410] <= 0.619863552;
cosLookup[9411] <= 0.619788312;
cosLookup[9412] <= 0.619713066;
cosLookup[9413] <= 0.619637814;
cosLookup[9414] <= 0.619562556;
cosLookup[9415] <= 0.619487293;
cosLookup[9416] <= 0.619412024;
cosLookup[9417] <= 0.619336749;
cosLookup[9418] <= 0.619261469;
cosLookup[9419] <= 0.619186183;
cosLookup[9420] <= 0.619110891;
cosLookup[9421] <= 0.619035593;
cosLookup[9422] <= 0.61896029;
cosLookup[9423] <= 0.618884981;
cosLookup[9424] <= 0.618809667;
cosLookup[9425] <= 0.618734346;
cosLookup[9426] <= 0.618659021;
cosLookup[9427] <= 0.618583689;
cosLookup[9428] <= 0.618508352;
cosLookup[9429] <= 0.618433009;
cosLookup[9430] <= 0.61835766;
cosLookup[9431] <= 0.618282306;
cosLookup[9432] <= 0.618206946;
cosLookup[9433] <= 0.61813158;
cosLookup[9434] <= 0.618056208;
cosLookup[9435] <= 0.617980831;
cosLookup[9436] <= 0.617905449;
cosLookup[9437] <= 0.61783006;
cosLookup[9438] <= 0.617754666;
cosLookup[9439] <= 0.617679266;
cosLookup[9440] <= 0.617603861;
cosLookup[9441] <= 0.61752845;
cosLookup[9442] <= 0.617453033;
cosLookup[9443] <= 0.61737761;
cosLookup[9444] <= 0.617302182;
cosLookup[9445] <= 0.617226748;
cosLookup[9446] <= 0.617151309;
cosLookup[9447] <= 0.617075863;
cosLookup[9448] <= 0.617000413;
cosLookup[9449] <= 0.616924956;
cosLookup[9450] <= 0.616849494;
cosLookup[9451] <= 0.616774026;
cosLookup[9452] <= 0.616698552;
cosLookup[9453] <= 0.616623073;
cosLookup[9454] <= 0.616547588;
cosLookup[9455] <= 0.616472098;
cosLookup[9456] <= 0.616396601;
cosLookup[9457] <= 0.616321099;
cosLookup[9458] <= 0.616245592;
cosLookup[9459] <= 0.616170079;
cosLookup[9460] <= 0.61609456;
cosLookup[9461] <= 0.616019035;
cosLookup[9462] <= 0.615943505;
cosLookup[9463] <= 0.615867969;
cosLookup[9464] <= 0.615792427;
cosLookup[9465] <= 0.61571688;
cosLookup[9466] <= 0.615641327;
cosLookup[9467] <= 0.615565769;
cosLookup[9468] <= 0.615490205;
cosLookup[9469] <= 0.615414635;
cosLookup[9470] <= 0.615339059;
cosLookup[9471] <= 0.615263478;
cosLookup[9472] <= 0.615187891;
cosLookup[9473] <= 0.615112299;
cosLookup[9474] <= 0.615036701;
cosLookup[9475] <= 0.614961097;
cosLookup[9476] <= 0.614885487;
cosLookup[9477] <= 0.614809872;
cosLookup[9478] <= 0.614734252;
cosLookup[9479] <= 0.614658625;
cosLookup[9480] <= 0.614582993;
cosLookup[9481] <= 0.614507355;
cosLookup[9482] <= 0.614431712;
cosLookup[9483] <= 0.614356063;
cosLookup[9484] <= 0.614280408;
cosLookup[9485] <= 0.614204748;
cosLookup[9486] <= 0.614129082;
cosLookup[9487] <= 0.614053411;
cosLookup[9488] <= 0.613977733;
cosLookup[9489] <= 0.613902051;
cosLookup[9490] <= 0.613826362;
cosLookup[9491] <= 0.613750668;
cosLookup[9492] <= 0.613674968;
cosLookup[9493] <= 0.613599263;
cosLookup[9494] <= 0.613523552;
cosLookup[9495] <= 0.613447835;
cosLookup[9496] <= 0.613372113;
cosLookup[9497] <= 0.613296385;
cosLookup[9498] <= 0.613220651;
cosLookup[9499] <= 0.613144912;
cosLookup[9500] <= 0.613069167;
cosLookup[9501] <= 0.612993416;
cosLookup[9502] <= 0.61291766;
cosLookup[9503] <= 0.612841898;
cosLookup[9504] <= 0.612766131;
cosLookup[9505] <= 0.612690358;
cosLookup[9506] <= 0.612614579;
cosLookup[9507] <= 0.612538795;
cosLookup[9508] <= 0.612463005;
cosLookup[9509] <= 0.612387209;
cosLookup[9510] <= 0.612311408;
cosLookup[9511] <= 0.612235601;
cosLookup[9512] <= 0.612159788;
cosLookup[9513] <= 0.61208397;
cosLookup[9514] <= 0.612008147;
cosLookup[9515] <= 0.611932317;
cosLookup[9516] <= 0.611856482;
cosLookup[9517] <= 0.611780642;
cosLookup[9518] <= 0.611704795;
cosLookup[9519] <= 0.611628943;
cosLookup[9520] <= 0.611553086;
cosLookup[9521] <= 0.611477223;
cosLookup[9522] <= 0.611401354;
cosLookup[9523] <= 0.61132548;
cosLookup[9524] <= 0.6112496;
cosLookup[9525] <= 0.611173714;
cosLookup[9526] <= 0.611097823;
cosLookup[9527] <= 0.611021926;
cosLookup[9528] <= 0.610946024;
cosLookup[9529] <= 0.610870116;
cosLookup[9530] <= 0.610794202;
cosLookup[9531] <= 0.610718283;
cosLookup[9532] <= 0.610642358;
cosLookup[9533] <= 0.610566427;
cosLookup[9534] <= 0.610490491;
cosLookup[9535] <= 0.610414549;
cosLookup[9536] <= 0.610338602;
cosLookup[9537] <= 0.610262649;
cosLookup[9538] <= 0.61018669;
cosLookup[9539] <= 0.610110726;
cosLookup[9540] <= 0.610034756;
cosLookup[9541] <= 0.609958781;
cosLookup[9542] <= 0.6098828;
cosLookup[9543] <= 0.609806813;
cosLookup[9544] <= 0.609730821;
cosLookup[9545] <= 0.609654823;
cosLookup[9546] <= 0.60957882;
cosLookup[9547] <= 0.609502811;
cosLookup[9548] <= 0.609426796;
cosLookup[9549] <= 0.609350776;
cosLookup[9550] <= 0.60927475;
cosLookup[9551] <= 0.609198719;
cosLookup[9552] <= 0.609122681;
cosLookup[9553] <= 0.609046639;
cosLookup[9554] <= 0.608970591;
cosLookup[9555] <= 0.608894537;
cosLookup[9556] <= 0.608818477;
cosLookup[9557] <= 0.608742412;
cosLookup[9558] <= 0.608666342;
cosLookup[9559] <= 0.608590265;
cosLookup[9560] <= 0.608514184;
cosLookup[9561] <= 0.608438096;
cosLookup[9562] <= 0.608362003;
cosLookup[9563] <= 0.608285904;
cosLookup[9564] <= 0.6082098;
cosLookup[9565] <= 0.60813369;
cosLookup[9566] <= 0.608057575;
cosLookup[9567] <= 0.607981454;
cosLookup[9568] <= 0.607905328;
cosLookup[9569] <= 0.607829195;
cosLookup[9570] <= 0.607753058;
cosLookup[9571] <= 0.607676914;
cosLookup[9572] <= 0.607600765;
cosLookup[9573] <= 0.607524611;
cosLookup[9574] <= 0.607448451;
cosLookup[9575] <= 0.607372285;
cosLookup[9576] <= 0.607296114;
cosLookup[9577] <= 0.607219937;
cosLookup[9578] <= 0.607143755;
cosLookup[9579] <= 0.607067567;
cosLookup[9580] <= 0.606991373;
cosLookup[9581] <= 0.606915174;
cosLookup[9582] <= 0.606838969;
cosLookup[9583] <= 0.606762759;
cosLookup[9584] <= 0.606686543;
cosLookup[9585] <= 0.606610322;
cosLookup[9586] <= 0.606534095;
cosLookup[9587] <= 0.606457862;
cosLookup[9588] <= 0.606381624;
cosLookup[9589] <= 0.60630538;
cosLookup[9590] <= 0.606229131;
cosLookup[9591] <= 0.606152876;
cosLookup[9592] <= 0.606076615;
cosLookup[9593] <= 0.606000349;
cosLookup[9594] <= 0.605924077;
cosLookup[9595] <= 0.6058478;
cosLookup[9596] <= 0.605771518;
cosLookup[9597] <= 0.605695229;
cosLookup[9598] <= 0.605618935;
cosLookup[9599] <= 0.605542636;
cosLookup[9600] <= 0.605466331;
cosLookup[9601] <= 0.60539002;
cosLookup[9602] <= 0.605313704;
cosLookup[9603] <= 0.605237382;
cosLookup[9604] <= 0.605161055;
cosLookup[9605] <= 0.605084722;
cosLookup[9606] <= 0.605008384;
cosLookup[9607] <= 0.60493204;
cosLookup[9608] <= 0.60485569;
cosLookup[9609] <= 0.604779335;
cosLookup[9610] <= 0.604702974;
cosLookup[9611] <= 0.604626608;
cosLookup[9612] <= 0.604550236;
cosLookup[9613] <= 0.604473859;
cosLookup[9614] <= 0.604397476;
cosLookup[9615] <= 0.604321088;
cosLookup[9616] <= 0.604244694;
cosLookup[9617] <= 0.604168294;
cosLookup[9618] <= 0.604091889;
cosLookup[9619] <= 0.604015478;
cosLookup[9620] <= 0.603939062;
cosLookup[9621] <= 0.60386264;
cosLookup[9622] <= 0.603786213;
cosLookup[9623] <= 0.60370978;
cosLookup[9624] <= 0.603633342;
cosLookup[9625] <= 0.603556898;
cosLookup[9626] <= 0.603480448;
cosLookup[9627] <= 0.603403993;
cosLookup[9628] <= 0.603327532;
cosLookup[9629] <= 0.603251066;
cosLookup[9630] <= 0.603174594;
cosLookup[9631] <= 0.603098117;
cosLookup[9632] <= 0.603021634;
cosLookup[9633] <= 0.602945146;
cosLookup[9634] <= 0.602868652;
cosLookup[9635] <= 0.602792153;
cosLookup[9636] <= 0.602715648;
cosLookup[9637] <= 0.602639137;
cosLookup[9638] <= 0.602562621;
cosLookup[9639] <= 0.6024861;
cosLookup[9640] <= 0.602409572;
cosLookup[9641] <= 0.60233304;
cosLookup[9642] <= 0.602256501;
cosLookup[9643] <= 0.602179958;
cosLookup[9644] <= 0.602103408;
cosLookup[9645] <= 0.602026854;
cosLookup[9646] <= 0.601950293;
cosLookup[9647] <= 0.601873727;
cosLookup[9648] <= 0.601797156;
cosLookup[9649] <= 0.601720579;
cosLookup[9650] <= 0.601643997;
cosLookup[9651] <= 0.601567409;
cosLookup[9652] <= 0.601490815;
cosLookup[9653] <= 0.601414216;
cosLookup[9654] <= 0.601337611;
cosLookup[9655] <= 0.601261001;
cosLookup[9656] <= 0.601184386;
cosLookup[9657] <= 0.601107764;
cosLookup[9658] <= 0.601031138;
cosLookup[9659] <= 0.600954505;
cosLookup[9660] <= 0.600877868;
cosLookup[9661] <= 0.600801224;
cosLookup[9662] <= 0.600724576;
cosLookup[9663] <= 0.600647921;
cosLookup[9664] <= 0.600571261;
cosLookup[9665] <= 0.600494596;
cosLookup[9666] <= 0.600417925;
cosLookup[9667] <= 0.600341249;
cosLookup[9668] <= 0.600264567;
cosLookup[9669] <= 0.600187879;
cosLookup[9670] <= 0.600111186;
cosLookup[9671] <= 0.600034488;
cosLookup[9672] <= 0.599957784;
cosLookup[9673] <= 0.599881074;
cosLookup[9674] <= 0.599804359;
cosLookup[9675] <= 0.599727639;
cosLookup[9676] <= 0.599650913;
cosLookup[9677] <= 0.599574181;
cosLookup[9678] <= 0.599497444;
cosLookup[9679] <= 0.599420701;
cosLookup[9680] <= 0.599343953;
cosLookup[9681] <= 0.5992672;
cosLookup[9682] <= 0.599190441;
cosLookup[9683] <= 0.599113676;
cosLookup[9684] <= 0.599036906;
cosLookup[9685] <= 0.59896013;
cosLookup[9686] <= 0.598883349;
cosLookup[9687] <= 0.598806562;
cosLookup[9688] <= 0.59872977;
cosLookup[9689] <= 0.598652973;
cosLookup[9690] <= 0.598576169;
cosLookup[9691] <= 0.598499361;
cosLookup[9692] <= 0.598422547;
cosLookup[9693] <= 0.598345727;
cosLookup[9694] <= 0.598268902;
cosLookup[9695] <= 0.598192071;
cosLookup[9696] <= 0.598115235;
cosLookup[9697] <= 0.598038393;
cosLookup[9698] <= 0.597961546;
cosLookup[9699] <= 0.597884693;
cosLookup[9700] <= 0.597807835;
cosLookup[9701] <= 0.597730972;
cosLookup[9702] <= 0.597654102;
cosLookup[9703] <= 0.597577228;
cosLookup[9704] <= 0.597500348;
cosLookup[9705] <= 0.597423462;
cosLookup[9706] <= 0.597346571;
cosLookup[9707] <= 0.597269674;
cosLookup[9708] <= 0.597192772;
cosLookup[9709] <= 0.597115865;
cosLookup[9710] <= 0.597038951;
cosLookup[9711] <= 0.596962033;
cosLookup[9712] <= 0.596885109;
cosLookup[9713] <= 0.596808179;
cosLookup[9714] <= 0.596731244;
cosLookup[9715] <= 0.596654304;
cosLookup[9716] <= 0.596577358;
cosLookup[9717] <= 0.596500406;
cosLookup[9718] <= 0.596423449;
cosLookup[9719] <= 0.596346487;
cosLookup[9720] <= 0.596269519;
cosLookup[9721] <= 0.596192545;
cosLookup[9722] <= 0.596115567;
cosLookup[9723] <= 0.596038582;
cosLookup[9724] <= 0.595961592;
cosLookup[9725] <= 0.595884597;
cosLookup[9726] <= 0.595807596;
cosLookup[9727] <= 0.59573059;
cosLookup[9728] <= 0.595653578;
cosLookup[9729] <= 0.595576561;
cosLookup[9730] <= 0.595499538;
cosLookup[9731] <= 0.59542251;
cosLookup[9732] <= 0.595345476;
cosLookup[9733] <= 0.595268437;
cosLookup[9734] <= 0.595191392;
cosLookup[9735] <= 0.595114342;
cosLookup[9736] <= 0.595037287;
cosLookup[9737] <= 0.594960226;
cosLookup[9738] <= 0.594883159;
cosLookup[9739] <= 0.594806087;
cosLookup[9740] <= 0.59472901;
cosLookup[9741] <= 0.594651927;
cosLookup[9742] <= 0.594574839;
cosLookup[9743] <= 0.594497745;
cosLookup[9744] <= 0.594420646;
cosLookup[9745] <= 0.594343541;
cosLookup[9746] <= 0.594266431;
cosLookup[9747] <= 0.594189315;
cosLookup[9748] <= 0.594112194;
cosLookup[9749] <= 0.594035067;
cosLookup[9750] <= 0.593957935;
cosLookup[9751] <= 0.593880797;
cosLookup[9752] <= 0.593803654;
cosLookup[9753] <= 0.593726506;
cosLookup[9754] <= 0.593649352;
cosLookup[9755] <= 0.593572193;
cosLookup[9756] <= 0.593495028;
cosLookup[9757] <= 0.593417858;
cosLookup[9758] <= 0.593340682;
cosLookup[9759] <= 0.593263501;
cosLookup[9760] <= 0.593186314;
cosLookup[9761] <= 0.593109122;
cosLookup[9762] <= 0.593031924;
cosLookup[9763] <= 0.592954721;
cosLookup[9764] <= 0.592877513;
cosLookup[9765] <= 0.592800299;
cosLookup[9766] <= 0.59272308;
cosLookup[9767] <= 0.592645855;
cosLookup[9768] <= 0.592568625;
cosLookup[9769] <= 0.592491389;
cosLookup[9770] <= 0.592414148;
cosLookup[9771] <= 0.592336901;
cosLookup[9772] <= 0.592259649;
cosLookup[9773] <= 0.592182392;
cosLookup[9774] <= 0.592105129;
cosLookup[9775] <= 0.59202786;
cosLookup[9776] <= 0.591950587;
cosLookup[9777] <= 0.591873307;
cosLookup[9778] <= 0.591796023;
cosLookup[9779] <= 0.591718733;
cosLookup[9780] <= 0.591641437;
cosLookup[9781] <= 0.591564136;
cosLookup[9782] <= 0.591486829;
cosLookup[9783] <= 0.591409518;
cosLookup[9784] <= 0.5913322;
cosLookup[9785] <= 0.591254878;
cosLookup[9786] <= 0.591177549;
cosLookup[9787] <= 0.591100216;
cosLookup[9788] <= 0.591022877;
cosLookup[9789] <= 0.590945532;
cosLookup[9790] <= 0.590868182;
cosLookup[9791] <= 0.590790827;
cosLookup[9792] <= 0.590713466;
cosLookup[9793] <= 0.5906361;
cosLookup[9794] <= 0.590558728;
cosLookup[9795] <= 0.590481351;
cosLookup[9796] <= 0.590403969;
cosLookup[9797] <= 0.590326581;
cosLookup[9798] <= 0.590249187;
cosLookup[9799] <= 0.590171788;
cosLookup[9800] <= 0.590094384;
cosLookup[9801] <= 0.590016975;
cosLookup[9802] <= 0.58993956;
cosLookup[9803] <= 0.589862139;
cosLookup[9804] <= 0.589784713;
cosLookup[9805] <= 0.589707282;
cosLookup[9806] <= 0.589629845;
cosLookup[9807] <= 0.589552403;
cosLookup[9808] <= 0.589474955;
cosLookup[9809] <= 0.589397502;
cosLookup[9810] <= 0.589320044;
cosLookup[9811] <= 0.58924258;
cosLookup[9812] <= 0.589165111;
cosLookup[9813] <= 0.589087636;
cosLookup[9814] <= 0.589010156;
cosLookup[9815] <= 0.58893267;
cosLookup[9816] <= 0.58885518;
cosLookup[9817] <= 0.588777683;
cosLookup[9818] <= 0.588700181;
cosLookup[9819] <= 0.588622674;
cosLookup[9820] <= 0.588545162;
cosLookup[9821] <= 0.588467644;
cosLookup[9822] <= 0.58839012;
cosLookup[9823] <= 0.588312592;
cosLookup[9824] <= 0.588235057;
cosLookup[9825] <= 0.588157518;
cosLookup[9826] <= 0.588079973;
cosLookup[9827] <= 0.588002422;
cosLookup[9828] <= 0.587924866;
cosLookup[9829] <= 0.587847305;
cosLookup[9830] <= 0.587769739;
cosLookup[9831] <= 0.587692166;
cosLookup[9832] <= 0.587614589;
cosLookup[9833] <= 0.587537006;
cosLookup[9834] <= 0.587459418;
cosLookup[9835] <= 0.587381824;
cosLookup[9836] <= 0.587304225;
cosLookup[9837] <= 0.587226621;
cosLookup[9838] <= 0.587149011;
cosLookup[9839] <= 0.587071396;
cosLookup[9840] <= 0.586993775;
cosLookup[9841] <= 0.586916149;
cosLookup[9842] <= 0.586838518;
cosLookup[9843] <= 0.586760881;
cosLookup[9844] <= 0.586683238;
cosLookup[9845] <= 0.586605591;
cosLookup[9846] <= 0.586527938;
cosLookup[9847] <= 0.586450279;
cosLookup[9848] <= 0.586372616;
cosLookup[9849] <= 0.586294946;
cosLookup[9850] <= 0.586217272;
cosLookup[9851] <= 0.586139592;
cosLookup[9852] <= 0.586061907;
cosLookup[9853] <= 0.585984216;
cosLookup[9854] <= 0.58590652;
cosLookup[9855] <= 0.585828818;
cosLookup[9856] <= 0.585751111;
cosLookup[9857] <= 0.585673399;
cosLookup[9858] <= 0.585595681;
cosLookup[9859] <= 0.585517958;
cosLookup[9860] <= 0.58544023;
cosLookup[9861] <= 0.585362496;
cosLookup[9862] <= 0.585284757;
cosLookup[9863] <= 0.585207012;
cosLookup[9864] <= 0.585129262;
cosLookup[9865] <= 0.585051507;
cosLookup[9866] <= 0.584973746;
cosLookup[9867] <= 0.58489598;
cosLookup[9868] <= 0.584818209;
cosLookup[9869] <= 0.584740432;
cosLookup[9870] <= 0.58466265;
cosLookup[9871] <= 0.584584862;
cosLookup[9872] <= 0.584507069;
cosLookup[9873] <= 0.584429271;
cosLookup[9874] <= 0.584351467;
cosLookup[9875] <= 0.584273658;
cosLookup[9876] <= 0.584195843;
cosLookup[9877] <= 0.584118024;
cosLookup[9878] <= 0.584040198;
cosLookup[9879] <= 0.583962368;
cosLookup[9880] <= 0.583884532;
cosLookup[9881] <= 0.583806691;
cosLookup[9882] <= 0.583728844;
cosLookup[9883] <= 0.583650992;
cosLookup[9884] <= 0.583573134;
cosLookup[9885] <= 0.583495272;
cosLookup[9886] <= 0.583417404;
cosLookup[9887] <= 0.58333953;
cosLookup[9888] <= 0.583261651;
cosLookup[9889] <= 0.583183767;
cosLookup[9890] <= 0.583105877;
cosLookup[9891] <= 0.583027982;
cosLookup[9892] <= 0.582950082;
cosLookup[9893] <= 0.582872176;
cosLookup[9894] <= 0.582794265;
cosLookup[9895] <= 0.582716349;
cosLookup[9896] <= 0.582638427;
cosLookup[9897] <= 0.5825605;
cosLookup[9898] <= 0.582482568;
cosLookup[9899] <= 0.58240463;
cosLookup[9900] <= 0.582326687;
cosLookup[9901] <= 0.582248738;
cosLookup[9902] <= 0.582170785;
cosLookup[9903] <= 0.582092825;
cosLookup[9904] <= 0.582014861;
cosLookup[9905] <= 0.581936891;
cosLookup[9906] <= 0.581858916;
cosLookup[9907] <= 0.581780935;
cosLookup[9908] <= 0.581702949;
cosLookup[9909] <= 0.581624958;
cosLookup[9910] <= 0.581546961;
cosLookup[9911] <= 0.581468959;
cosLookup[9912] <= 0.581390952;
cosLookup[9913] <= 0.581312939;
cosLookup[9914] <= 0.581234921;
cosLookup[9915] <= 0.581156898;
cosLookup[9916] <= 0.581078869;
cosLookup[9917] <= 0.581000835;
cosLookup[9918] <= 0.580922795;
cosLookup[9919] <= 0.580844751;
cosLookup[9920] <= 0.580766701;
cosLookup[9921] <= 0.580688645;
cosLookup[9922] <= 0.580610584;
cosLookup[9923] <= 0.580532518;
cosLookup[9924] <= 0.580454447;
cosLookup[9925] <= 0.58037637;
cosLookup[9926] <= 0.580298288;
cosLookup[9927] <= 0.580220201;
cosLookup[9928] <= 0.580142108;
cosLookup[9929] <= 0.58006401;
cosLookup[9930] <= 0.579985906;
cosLookup[9931] <= 0.579907797;
cosLookup[9932] <= 0.579829683;
cosLookup[9933] <= 0.579751564;
cosLookup[9934] <= 0.579673439;
cosLookup[9935] <= 0.579595309;
cosLookup[9936] <= 0.579517174;
cosLookup[9937] <= 0.579439033;
cosLookup[9938] <= 0.579360887;
cosLookup[9939] <= 0.579282735;
cosLookup[9940] <= 0.579204579;
cosLookup[9941] <= 0.579126417;
cosLookup[9942] <= 0.579048249;
cosLookup[9943] <= 0.578970077;
cosLookup[9944] <= 0.578891899;
cosLookup[9945] <= 0.578813715;
cosLookup[9946] <= 0.578735527;
cosLookup[9947] <= 0.578657333;
cosLookup[9948] <= 0.578579133;
cosLookup[9949] <= 0.578500929;
cosLookup[9950] <= 0.578422719;
cosLookup[9951] <= 0.578344503;
cosLookup[9952] <= 0.578266283;
cosLookup[9953] <= 0.578188057;
cosLookup[9954] <= 0.578109826;
cosLookup[9955] <= 0.578031589;
cosLookup[9956] <= 0.577953347;
cosLookup[9957] <= 0.5778751;
cosLookup[9958] <= 0.577796848;
cosLookup[9959] <= 0.57771859;
cosLookup[9960] <= 0.577640327;
cosLookup[9961] <= 0.577562059;
cosLookup[9962] <= 0.577483785;
cosLookup[9963] <= 0.577405506;
cosLookup[9964] <= 0.577327222;
cosLookup[9965] <= 0.577248932;
cosLookup[9966] <= 0.577170637;
cosLookup[9967] <= 0.577092337;
cosLookup[9968] <= 0.577014031;
cosLookup[9969] <= 0.57693572;
cosLookup[9970] <= 0.576857404;
cosLookup[9971] <= 0.576779083;
cosLookup[9972] <= 0.576700756;
cosLookup[9973] <= 0.576622424;
cosLookup[9974] <= 0.576544087;
cosLookup[9975] <= 0.576465744;
cosLookup[9976] <= 0.576387396;
cosLookup[9977] <= 0.576309043;
cosLookup[9978] <= 0.576230684;
cosLookup[9979] <= 0.57615232;
cosLookup[9980] <= 0.576073951;
cosLookup[9981] <= 0.575995577;
cosLookup[9982] <= 0.575917197;
cosLookup[9983] <= 0.575838812;
cosLookup[9984] <= 0.575760422;
cosLookup[9985] <= 0.575682026;
cosLookup[9986] <= 0.575603625;
cosLookup[9987] <= 0.575525219;
cosLookup[9988] <= 0.575446807;
cosLookup[9989] <= 0.575368391;
cosLookup[9990] <= 0.575289969;
cosLookup[9991] <= 0.575211541;
cosLookup[9992] <= 0.575133109;
cosLookup[9993] <= 0.575054671;
cosLookup[9994] <= 0.574976227;
cosLookup[9995] <= 0.574897779;
cosLookup[9996] <= 0.574819325;
cosLookup[9997] <= 0.574740866;
cosLookup[9998] <= 0.574662402;
cosLookup[9999] <= 0.574583932;
cosLookup[10000] <= 0.574505457;
cosLookup[10001] <= 0.574426977;
cosLookup[10002] <= 0.574348491;
cosLookup[10003] <= 0.574270001;
cosLookup[10004] <= 0.574191505;
cosLookup[10005] <= 0.574113003;
cosLookup[10006] <= 0.574034497;
cosLookup[10007] <= 0.573955985;
cosLookup[10008] <= 0.573877468;
cosLookup[10009] <= 0.573798945;
cosLookup[10010] <= 0.573720418;
cosLookup[10011] <= 0.573641885;
cosLookup[10012] <= 0.573563346;
cosLookup[10013] <= 0.573484803;
cosLookup[10014] <= 0.573406254;
cosLookup[10015] <= 0.5733277;
cosLookup[10016] <= 0.573249141;
cosLookup[10017] <= 0.573170576;
cosLookup[10018] <= 0.573092006;
cosLookup[10019] <= 0.573013431;
cosLookup[10020] <= 0.57293485;
cosLookup[10021] <= 0.572856265;
cosLookup[10022] <= 0.572777674;
cosLookup[10023] <= 0.572699078;
cosLookup[10024] <= 0.572620476;
cosLookup[10025] <= 0.572541869;
cosLookup[10026] <= 0.572463257;
cosLookup[10027] <= 0.57238464;
cosLookup[10028] <= 0.572306018;
cosLookup[10029] <= 0.57222739;
cosLookup[10030] <= 0.572148757;
cosLookup[10031] <= 0.572070118;
cosLookup[10032] <= 0.571991475;
cosLookup[10033] <= 0.571912826;
cosLookup[10034] <= 0.571834172;
cosLookup[10035] <= 0.571755513;
cosLookup[10036] <= 0.571676848;
cosLookup[10037] <= 0.571598178;
cosLookup[10038] <= 0.571519503;
cosLookup[10039] <= 0.571440823;
cosLookup[10040] <= 0.571362137;
cosLookup[10041] <= 0.571283446;
cosLookup[10042] <= 0.57120475;
cosLookup[10043] <= 0.571126049;
cosLookup[10044] <= 0.571047342;
cosLookup[10045] <= 0.57096863;
cosLookup[10046] <= 0.570889913;
cosLookup[10047] <= 0.570811191;
cosLookup[10048] <= 0.570732463;
cosLookup[10049] <= 0.57065373;
cosLookup[10050] <= 0.570574992;
cosLookup[10051] <= 0.570496249;
cosLookup[10052] <= 0.5704175;
cosLookup[10053] <= 0.570338746;
cosLookup[10054] <= 0.570259987;
cosLookup[10055] <= 0.570181223;
cosLookup[10056] <= 0.570102453;
cosLookup[10057] <= 0.570023679;
cosLookup[10058] <= 0.569944898;
cosLookup[10059] <= 0.569866113;
cosLookup[10060] <= 0.569787323;
cosLookup[10061] <= 0.569708527;
cosLookup[10062] <= 0.569629726;
cosLookup[10063] <= 0.56955092;
cosLookup[10064] <= 0.569472108;
cosLookup[10065] <= 0.569393291;
cosLookup[10066] <= 0.56931447;
cosLookup[10067] <= 0.569235642;
cosLookup[10068] <= 0.56915681;
cosLookup[10069] <= 0.569077972;
cosLookup[10070] <= 0.568999129;
cosLookup[10071] <= 0.568920281;
cosLookup[10072] <= 0.568841428;
cosLookup[10073] <= 0.568762569;
cosLookup[10074] <= 0.568683706;
cosLookup[10075] <= 0.568604837;
cosLookup[10076] <= 0.568525962;
cosLookup[10077] <= 0.568447083;
cosLookup[10078] <= 0.568368198;
cosLookup[10079] <= 0.568289308;
cosLookup[10080] <= 0.568210413;
cosLookup[10081] <= 0.568131513;
cosLookup[10082] <= 0.568052607;
cosLookup[10083] <= 0.567973696;
cosLookup[10084] <= 0.56789478;
cosLookup[10085] <= 0.567815859;
cosLookup[10086] <= 0.567736932;
cosLookup[10087] <= 0.567658001;
cosLookup[10088] <= 0.567579064;
cosLookup[10089] <= 0.567500122;
cosLookup[10090] <= 0.567421174;
cosLookup[10091] <= 0.567342222;
cosLookup[10092] <= 0.567263264;
cosLookup[10093] <= 0.567184301;
cosLookup[10094] <= 0.567105333;
cosLookup[10095] <= 0.567026359;
cosLookup[10096] <= 0.566947381;
cosLookup[10097] <= 0.566868397;
cosLookup[10098] <= 0.566789408;
cosLookup[10099] <= 0.566710414;
cosLookup[10100] <= 0.566631414;
cosLookup[10101] <= 0.566552409;
cosLookup[10102] <= 0.566473399;
cosLookup[10103] <= 0.566394384;
cosLookup[10104] <= 0.566315364;
cosLookup[10105] <= 0.566236338;
cosLookup[10106] <= 0.566157308;
cosLookup[10107] <= 0.566078272;
cosLookup[10108] <= 0.565999231;
cosLookup[10109] <= 0.565920184;
cosLookup[10110] <= 0.565841133;
cosLookup[10111] <= 0.565762076;
cosLookup[10112] <= 0.565683014;
cosLookup[10113] <= 0.565603947;
cosLookup[10114] <= 0.565524875;
cosLookup[10115] <= 0.565445797;
cosLookup[10116] <= 0.565366714;
cosLookup[10117] <= 0.565287626;
cosLookup[10118] <= 0.565208533;
cosLookup[10119] <= 0.565129435;
cosLookup[10120] <= 0.565050331;
cosLookup[10121] <= 0.564971223;
cosLookup[10122] <= 0.564892109;
cosLookup[10123] <= 0.56481299;
cosLookup[10124] <= 0.564733865;
cosLookup[10125] <= 0.564654736;
cosLookup[10126] <= 0.564575601;
cosLookup[10127] <= 0.564496461;
cosLookup[10128] <= 0.564417316;
cosLookup[10129] <= 0.564338166;
cosLookup[10130] <= 0.564259011;
cosLookup[10131] <= 0.56417985;
cosLookup[10132] <= 0.564100684;
cosLookup[10133] <= 0.564021513;
cosLookup[10134] <= 0.563942337;
cosLookup[10135] <= 0.563863156;
cosLookup[10136] <= 0.563783969;
cosLookup[10137] <= 0.563704777;
cosLookup[10138] <= 0.56362558;
cosLookup[10139] <= 0.563546378;
cosLookup[10140] <= 0.563467171;
cosLookup[10141] <= 0.563387959;
cosLookup[10142] <= 0.563308741;
cosLookup[10143] <= 0.563229518;
cosLookup[10144] <= 0.56315029;
cosLookup[10145] <= 0.563071057;
cosLookup[10146] <= 0.562991819;
cosLookup[10147] <= 0.562912575;
cosLookup[10148] <= 0.562833326;
cosLookup[10149] <= 0.562754073;
cosLookup[10150] <= 0.562674813;
cosLookup[10151] <= 0.562595549;
cosLookup[10152] <= 0.56251628;
cosLookup[10153] <= 0.562437005;
cosLookup[10154] <= 0.562357726;
cosLookup[10155] <= 0.562278441;
cosLookup[10156] <= 0.562199151;
cosLookup[10157] <= 0.562119855;
cosLookup[10158] <= 0.562040555;
cosLookup[10159] <= 0.561961249;
cosLookup[10160] <= 0.561881939;
cosLookup[10161] <= 0.561802623;
cosLookup[10162] <= 0.561723302;
cosLookup[10163] <= 0.561643975;
cosLookup[10164] <= 0.561564644;
cosLookup[10165] <= 0.561485308;
cosLookup[10166] <= 0.561405966;
cosLookup[10167] <= 0.561326619;
cosLookup[10168] <= 0.561247267;
cosLookup[10169] <= 0.56116791;
cosLookup[10170] <= 0.561088547;
cosLookup[10171] <= 0.56100918;
cosLookup[10172] <= 0.560929807;
cosLookup[10173] <= 0.560850429;
cosLookup[10174] <= 0.560771046;
cosLookup[10175] <= 0.560691658;
cosLookup[10176] <= 0.560612265;
cosLookup[10177] <= 0.560532866;
cosLookup[10178] <= 0.560453463;
cosLookup[10179] <= 0.560374054;
cosLookup[10180] <= 0.56029464;
cosLookup[10181] <= 0.560215221;
cosLookup[10182] <= 0.560135797;
cosLookup[10183] <= 0.560056368;
cosLookup[10184] <= 0.559976933;
cosLookup[10185] <= 0.559897493;
cosLookup[10186] <= 0.559818049;
cosLookup[10187] <= 0.559738599;
cosLookup[10188] <= 0.559659144;
cosLookup[10189] <= 0.559579683;
cosLookup[10190] <= 0.559500218;
cosLookup[10191] <= 0.559420747;
cosLookup[10192] <= 0.559341272;
cosLookup[10193] <= 0.559261791;
cosLookup[10194] <= 0.559182305;
cosLookup[10195] <= 0.559102814;
cosLookup[10196] <= 0.559023318;
cosLookup[10197] <= 0.558943816;
cosLookup[10198] <= 0.55886431;
cosLookup[10199] <= 0.558784798;
cosLookup[10200] <= 0.558705281;
cosLookup[10201] <= 0.55862576;
cosLookup[10202] <= 0.558546232;
cosLookup[10203] <= 0.5584667;
cosLookup[10204] <= 0.558387163;
cosLookup[10205] <= 0.558307621;
cosLookup[10206] <= 0.558228073;
cosLookup[10207] <= 0.55814852;
cosLookup[10208] <= 0.558068962;
cosLookup[10209] <= 0.557989399;
cosLookup[10210] <= 0.557909831;
cosLookup[10211] <= 0.557830258;
cosLookup[10212] <= 0.55775068;
cosLookup[10213] <= 0.557671096;
cosLookup[10214] <= 0.557591508;
cosLookup[10215] <= 0.557511914;
cosLookup[10216] <= 0.557432315;
cosLookup[10217] <= 0.557352711;
cosLookup[10218] <= 0.557273102;
cosLookup[10219] <= 0.557193488;
cosLookup[10220] <= 0.557113868;
cosLookup[10221] <= 0.557034244;
cosLookup[10222] <= 0.556954614;
cosLookup[10223] <= 0.556874979;
cosLookup[10224] <= 0.55679534;
cosLookup[10225] <= 0.556715695;
cosLookup[10226] <= 0.556636044;
cosLookup[10227] <= 0.556556389;
cosLookup[10228] <= 0.556476729;
cosLookup[10229] <= 0.556397064;
cosLookup[10230] <= 0.556317393;
cosLookup[10231] <= 0.556237717;
cosLookup[10232] <= 0.556158037;
cosLookup[10233] <= 0.556078351;
cosLookup[10234] <= 0.55599866;
cosLookup[10235] <= 0.555918964;
cosLookup[10236] <= 0.555839262;
cosLookup[10237] <= 0.555759556;
cosLookup[10238] <= 0.555679845;
cosLookup[10239] <= 0.555600128;
cosLookup[10240] <= 0.555520406;
cosLookup[10241] <= 0.55544068;
cosLookup[10242] <= 0.555360948;
cosLookup[10243] <= 0.555281211;
cosLookup[10244] <= 0.555201469;
cosLookup[10245] <= 0.555121722;
cosLookup[10246] <= 0.555041969;
cosLookup[10247] <= 0.554962212;
cosLookup[10248] <= 0.554882449;
cosLookup[10249] <= 0.554802682;
cosLookup[10250] <= 0.554722909;
cosLookup[10251] <= 0.554643131;
cosLookup[10252] <= 0.554563348;
cosLookup[10253] <= 0.55448356;
cosLookup[10254] <= 0.554403767;
cosLookup[10255] <= 0.554323969;
cosLookup[10256] <= 0.554244166;
cosLookup[10257] <= 0.554164358;
cosLookup[10258] <= 0.554084544;
cosLookup[10259] <= 0.554004725;
cosLookup[10260] <= 0.553924902;
cosLookup[10261] <= 0.553845073;
cosLookup[10262] <= 0.553765239;
cosLookup[10263] <= 0.5536854;
cosLookup[10264] <= 0.553605556;
cosLookup[10265] <= 0.553525707;
cosLookup[10266] <= 0.553445853;
cosLookup[10267] <= 0.553365994;
cosLookup[10268] <= 0.553286129;
cosLookup[10269] <= 0.55320626;
cosLookup[10270] <= 0.553126385;
cosLookup[10271] <= 0.553046506;
cosLookup[10272] <= 0.552966621;
cosLookup[10273] <= 0.552886731;
cosLookup[10274] <= 0.552806836;
cosLookup[10275] <= 0.552726936;
cosLookup[10276] <= 0.552647031;
cosLookup[10277] <= 0.552567121;
cosLookup[10278] <= 0.552487206;
cosLookup[10279] <= 0.552407286;
cosLookup[10280] <= 0.55232736;
cosLookup[10281] <= 0.55224743;
cosLookup[10282] <= 0.552167494;
cosLookup[10283] <= 0.552087554;
cosLookup[10284] <= 0.552007608;
cosLookup[10285] <= 0.551927657;
cosLookup[10286] <= 0.551847702;
cosLookup[10287] <= 0.551767741;
cosLookup[10288] <= 0.551687775;
cosLookup[10289] <= 0.551607804;
cosLookup[10290] <= 0.551527828;
cosLookup[10291] <= 0.551447847;
cosLookup[10292] <= 0.55136786;
cosLookup[10293] <= 0.551287869;
cosLookup[10294] <= 0.551207873;
cosLookup[10295] <= 0.551127871;
cosLookup[10296] <= 0.551047865;
cosLookup[10297] <= 0.550967853;
cosLookup[10298] <= 0.550887836;
cosLookup[10299] <= 0.550807815;
cosLookup[10300] <= 0.550727788;
cosLookup[10301] <= 0.550647756;
cosLookup[10302] <= 0.550567719;
cosLookup[10303] <= 0.550487677;
cosLookup[10304] <= 0.55040763;
cosLookup[10305] <= 0.550327578;
cosLookup[10306] <= 0.550247521;
cosLookup[10307] <= 0.550167459;
cosLookup[10308] <= 0.550087392;
cosLookup[10309] <= 0.550007319;
cosLookup[10310] <= 0.549927242;
cosLookup[10311] <= 0.54984716;
cosLookup[10312] <= 0.549767072;
cosLookup[10313] <= 0.54968698;
cosLookup[10314] <= 0.549606882;
cosLookup[10315] <= 0.549526779;
cosLookup[10316] <= 0.549446672;
cosLookup[10317] <= 0.549366559;
cosLookup[10318] <= 0.549286441;
cosLookup[10319] <= 0.549206318;
cosLookup[10320] <= 0.54912619;
cosLookup[10321] <= 0.549046057;
cosLookup[10322] <= 0.54896592;
cosLookup[10323] <= 0.548885776;
cosLookup[10324] <= 0.548805628;
cosLookup[10325] <= 0.548725475;
cosLookup[10326] <= 0.548645317;
cosLookup[10327] <= 0.548565154;
cosLookup[10328] <= 0.548484986;
cosLookup[10329] <= 0.548404812;
cosLookup[10330] <= 0.548324634;
cosLookup[10331] <= 0.548244451;
cosLookup[10332] <= 0.548164262;
cosLookup[10333] <= 0.548084069;
cosLookup[10334] <= 0.54800387;
cosLookup[10335] <= 0.547923667;
cosLookup[10336] <= 0.547843458;
cosLookup[10337] <= 0.547763245;
cosLookup[10338] <= 0.547683026;
cosLookup[10339] <= 0.547602802;
cosLookup[10340] <= 0.547522574;
cosLookup[10341] <= 0.54744234;
cosLookup[10342] <= 0.547362101;
cosLookup[10343] <= 0.547281857;
cosLookup[10344] <= 0.547201609;
cosLookup[10345] <= 0.547121355;
cosLookup[10346] <= 0.547041096;
cosLookup[10347] <= 0.546960832;
cosLookup[10348] <= 0.546880563;
cosLookup[10349] <= 0.546800289;
cosLookup[10350] <= 0.54672001;
cosLookup[10351] <= 0.546639726;
cosLookup[10352] <= 0.546559437;
cosLookup[10353] <= 0.546479143;
cosLookup[10354] <= 0.546398844;
cosLookup[10355] <= 0.54631854;
cosLookup[10356] <= 0.54623823;
cosLookup[10357] <= 0.546157916;
cosLookup[10358] <= 0.546077597;
cosLookup[10359] <= 0.545997273;
cosLookup[10360] <= 0.545916944;
cosLookup[10361] <= 0.545836609;
cosLookup[10362] <= 0.54575627;
cosLookup[10363] <= 0.545675926;
cosLookup[10364] <= 0.545595576;
cosLookup[10365] <= 0.545515222;
cosLookup[10366] <= 0.545434863;
cosLookup[10367] <= 0.545354498;
cosLookup[10368] <= 0.545274129;
cosLookup[10369] <= 0.545193755;
cosLookup[10370] <= 0.545113375;
cosLookup[10371] <= 0.545032991;
cosLookup[10372] <= 0.544952602;
cosLookup[10373] <= 0.544872207;
cosLookup[10374] <= 0.544791808;
cosLookup[10375] <= 0.544711403;
cosLookup[10376] <= 0.544630994;
cosLookup[10377] <= 0.544550579;
cosLookup[10378] <= 0.54447016;
cosLookup[10379] <= 0.544389735;
cosLookup[10380] <= 0.544309306;
cosLookup[10381] <= 0.544228872;
cosLookup[10382] <= 0.544148432;
cosLookup[10383] <= 0.544067988;
cosLookup[10384] <= 0.543987538;
cosLookup[10385] <= 0.543907084;
cosLookup[10386] <= 0.543826624;
cosLookup[10387] <= 0.54374616;
cosLookup[10388] <= 0.54366569;
cosLookup[10389] <= 0.543585216;
cosLookup[10390] <= 0.543504736;
cosLookup[10391] <= 0.543424252;
cosLookup[10392] <= 0.543343762;
cosLookup[10393] <= 0.543263268;
cosLookup[10394] <= 0.543182769;
cosLookup[10395] <= 0.543102264;
cosLookup[10396] <= 0.543021755;
cosLookup[10397] <= 0.54294124;
cosLookup[10398] <= 0.542860721;
cosLookup[10399] <= 0.542780196;
cosLookup[10400] <= 0.542699667;
cosLookup[10401] <= 0.542619133;
cosLookup[10402] <= 0.542538593;
cosLookup[10403] <= 0.542458049;
cosLookup[10404] <= 0.5423775;
cosLookup[10405] <= 0.542296945;
cosLookup[10406] <= 0.542216386;
cosLookup[10407] <= 0.542135822;
cosLookup[10408] <= 0.542055252;
cosLookup[10409] <= 0.541974678;
cosLookup[10410] <= 0.541894099;
cosLookup[10411] <= 0.541813515;
cosLookup[10412] <= 0.541732925;
cosLookup[10413] <= 0.541652331;
cosLookup[10414] <= 0.541571732;
cosLookup[10415] <= 0.541491128;
cosLookup[10416] <= 0.541410519;
cosLookup[10417] <= 0.541329905;
cosLookup[10418] <= 0.541249285;
cosLookup[10419] <= 0.541168661;
cosLookup[10420] <= 0.541088032;
cosLookup[10421] <= 0.541007398;
cosLookup[10422] <= 0.540926759;
cosLookup[10423] <= 0.540846115;
cosLookup[10424] <= 0.540765466;
cosLookup[10425] <= 0.540684813;
cosLookup[10426] <= 0.540604154;
cosLookup[10427] <= 0.54052349;
cosLookup[10428] <= 0.540442821;
cosLookup[10429] <= 0.540362147;
cosLookup[10430] <= 0.540281469;
cosLookup[10431] <= 0.540200785;
cosLookup[10432] <= 0.540120096;
cosLookup[10433] <= 0.540039403;
cosLookup[10434] <= 0.539958704;
cosLookup[10435] <= 0.539878;
cosLookup[10436] <= 0.539797292;
cosLookup[10437] <= 0.539716578;
cosLookup[10438] <= 0.53963586;
cosLookup[10439] <= 0.539555136;
cosLookup[10440] <= 0.539474408;
cosLookup[10441] <= 0.539393675;
cosLookup[10442] <= 0.539312936;
cosLookup[10443] <= 0.539232193;
cosLookup[10444] <= 0.539151445;
cosLookup[10445] <= 0.539070692;
cosLookup[10446] <= 0.538989934;
cosLookup[10447] <= 0.538909171;
cosLookup[10448] <= 0.538828403;
cosLookup[10449] <= 0.53874763;
cosLookup[10450] <= 0.538666852;
cosLookup[10451] <= 0.538586069;
cosLookup[10452] <= 0.538505281;
cosLookup[10453] <= 0.538424488;
cosLookup[10454] <= 0.53834369;
cosLookup[10455] <= 0.538262888;
cosLookup[10456] <= 0.53818208;
cosLookup[10457] <= 0.538101267;
cosLookup[10458] <= 0.53802045;
cosLookup[10459] <= 0.537939627;
cosLookup[10460] <= 0.5378588;
cosLookup[10461] <= 0.537777968;
cosLookup[10462] <= 0.53769713;
cosLookup[10463] <= 0.537616288;
cosLookup[10464] <= 0.537535441;
cosLookup[10465] <= 0.537454589;
cosLookup[10466] <= 0.537373732;
cosLookup[10467] <= 0.53729287;
cosLookup[10468] <= 0.537212003;
cosLookup[10469] <= 0.537131131;
cosLookup[10470] <= 0.537050254;
cosLookup[10471] <= 0.536969372;
cosLookup[10472] <= 0.536888485;
cosLookup[10473] <= 0.536807594;
cosLookup[10474] <= 0.536726697;
cosLookup[10475] <= 0.536645796;
cosLookup[10476] <= 0.536564889;
cosLookup[10477] <= 0.536483978;
cosLookup[10478] <= 0.536403062;
cosLookup[10479] <= 0.53632214;
cosLookup[10480] <= 0.536241214;
cosLookup[10481] <= 0.536160283;
cosLookup[10482] <= 0.536079347;
cosLookup[10483] <= 0.535998406;
cosLookup[10484] <= 0.53591746;
cosLookup[10485] <= 0.535836509;
cosLookup[10486] <= 0.535755554;
cosLookup[10487] <= 0.535674593;
cosLookup[10488] <= 0.535593627;
cosLookup[10489] <= 0.535512657;
cosLookup[10490] <= 0.535431681;
cosLookup[10491] <= 0.535350701;
cosLookup[10492] <= 0.535269716;
cosLookup[10493] <= 0.535188726;
cosLookup[10494] <= 0.535107731;
cosLookup[10495] <= 0.53502673;
cosLookup[10496] <= 0.534945726;
cosLookup[10497] <= 0.534864716;
cosLookup[10498] <= 0.534783701;
cosLookup[10499] <= 0.534702681;
cosLookup[10500] <= 0.534621657;
cosLookup[10501] <= 0.534540627;
cosLookup[10502] <= 0.534459593;
cosLookup[10503] <= 0.534378553;
cosLookup[10504] <= 0.534297509;
cosLookup[10505] <= 0.53421646;
cosLookup[10506] <= 0.534135406;
cosLookup[10507] <= 0.534054347;
cosLookup[10508] <= 0.533973283;
cosLookup[10509] <= 0.533892214;
cosLookup[10510] <= 0.53381114;
cosLookup[10511] <= 0.533730061;
cosLookup[10512] <= 0.533648978;
cosLookup[10513] <= 0.533567889;
cosLookup[10514] <= 0.533486796;
cosLookup[10515] <= 0.533405698;
cosLookup[10516] <= 0.533324595;
cosLookup[10517] <= 0.533243487;
cosLookup[10518] <= 0.533162374;
cosLookup[10519] <= 0.533081256;
cosLookup[10520] <= 0.533000133;
cosLookup[10521] <= 0.532919005;
cosLookup[10522] <= 0.532837873;
cosLookup[10523] <= 0.532756735;
cosLookup[10524] <= 0.532675593;
cosLookup[10525] <= 0.532594446;
cosLookup[10526] <= 0.532513293;
cosLookup[10527] <= 0.532432136;
cosLookup[10528] <= 0.532350974;
cosLookup[10529] <= 0.532269808;
cosLookup[10530] <= 0.532188636;
cosLookup[10531] <= 0.532107459;
cosLookup[10532] <= 0.532026278;
cosLookup[10533] <= 0.531945091;
cosLookup[10534] <= 0.5318639;
cosLookup[10535] <= 0.531782704;
cosLookup[10536] <= 0.531701503;
cosLookup[10537] <= 0.531620297;
cosLookup[10538] <= 0.531539086;
cosLookup[10539] <= 0.53145787;
cosLookup[10540] <= 0.531376649;
cosLookup[10541] <= 0.531295424;
cosLookup[10542] <= 0.531214194;
cosLookup[10543] <= 0.531132958;
cosLookup[10544] <= 0.531051718;
cosLookup[10545] <= 0.530970473;
cosLookup[10546] <= 0.530889223;
cosLookup[10547] <= 0.530807968;
cosLookup[10548] <= 0.530726709;
cosLookup[10549] <= 0.530645444;
cosLookup[10550] <= 0.530564175;
cosLookup[10551] <= 0.5304829;
cosLookup[10552] <= 0.530401621;
cosLookup[10553] <= 0.530320337;
cosLookup[10554] <= 0.530239048;
cosLookup[10555] <= 0.530157754;
cosLookup[10556] <= 0.530076456;
cosLookup[10557] <= 0.529995152;
cosLookup[10558] <= 0.529913844;
cosLookup[10559] <= 0.52983253;
cosLookup[10560] <= 0.529751212;
cosLookup[10561] <= 0.529669889;
cosLookup[10562] <= 0.529588561;
cosLookup[10563] <= 0.529507228;
cosLookup[10564] <= 0.529425891;
cosLookup[10565] <= 0.529344548;
cosLookup[10566] <= 0.529263201;
cosLookup[10567] <= 0.529181848;
cosLookup[10568] <= 0.529100491;
cosLookup[10569] <= 0.529019129;
cosLookup[10570] <= 0.528937762;
cosLookup[10571] <= 0.528856391;
cosLookup[10572] <= 0.528775014;
cosLookup[10573] <= 0.528693633;
cosLookup[10574] <= 0.528612246;
cosLookup[10575] <= 0.528530855;
cosLookup[10576] <= 0.528449459;
cosLookup[10577] <= 0.528368058;
cosLookup[10578] <= 0.528286653;
cosLookup[10579] <= 0.528205242;
cosLookup[10580] <= 0.528123827;
cosLookup[10581] <= 0.528042406;
cosLookup[10582] <= 0.527960981;
cosLookup[10583] <= 0.527879551;
cosLookup[10584] <= 0.527798116;
cosLookup[10585] <= 0.527716677;
cosLookup[10586] <= 0.527635232;
cosLookup[10587] <= 0.527553783;
cosLookup[10588] <= 0.527472328;
cosLookup[10589] <= 0.527390869;
cosLookup[10590] <= 0.527309405;
cosLookup[10591] <= 0.527227936;
cosLookup[10592] <= 0.527146463;
cosLookup[10593] <= 0.527064984;
cosLookup[10594] <= 0.526983501;
cosLookup[10595] <= 0.526902013;
cosLookup[10596] <= 0.52682052;
cosLookup[10597] <= 0.526739022;
cosLookup[10598] <= 0.526657519;
cosLookup[10599] <= 0.526576012;
cosLookup[10600] <= 0.526494499;
cosLookup[10601] <= 0.526412982;
cosLookup[10602] <= 0.52633146;
cosLookup[10603] <= 0.526249933;
cosLookup[10604] <= 0.526168401;
cosLookup[10605] <= 0.526086865;
cosLookup[10606] <= 0.526005323;
cosLookup[10607] <= 0.525923777;
cosLookup[10608] <= 0.525842226;
cosLookup[10609] <= 0.52576067;
cosLookup[10610] <= 0.525679109;
cosLookup[10611] <= 0.525597543;
cosLookup[10612] <= 0.525515973;
cosLookup[10613] <= 0.525434398;
cosLookup[10614] <= 0.525352818;
cosLookup[10615] <= 0.525271233;
cosLookup[10616] <= 0.525189643;
cosLookup[10617] <= 0.525108048;
cosLookup[10618] <= 0.525026449;
cosLookup[10619] <= 0.524944845;
cosLookup[10620] <= 0.524863236;
cosLookup[10621] <= 0.524781622;
cosLookup[10622] <= 0.524700003;
cosLookup[10623] <= 0.52461838;
cosLookup[10624] <= 0.524536751;
cosLookup[10625] <= 0.524455118;
cosLookup[10626] <= 0.52437348;
cosLookup[10627] <= 0.524291837;
cosLookup[10628] <= 0.52421019;
cosLookup[10629] <= 0.524128537;
cosLookup[10630] <= 0.52404688;
cosLookup[10631] <= 0.523965218;
cosLookup[10632] <= 0.523883551;
cosLookup[10633] <= 0.523801879;
cosLookup[10634] <= 0.523720203;
cosLookup[10635] <= 0.523638521;
cosLookup[10636] <= 0.523556835;
cosLookup[10637] <= 0.523475144;
cosLookup[10638] <= 0.523393448;
cosLookup[10639] <= 0.523311748;
cosLookup[10640] <= 0.523230042;
cosLookup[10641] <= 0.523148332;
cosLookup[10642] <= 0.523066617;
cosLookup[10643] <= 0.522984897;
cosLookup[10644] <= 0.522903173;
cosLookup[10645] <= 0.522821443;
cosLookup[10646] <= 0.522739709;
cosLookup[10647] <= 0.52265797;
cosLookup[10648] <= 0.522576226;
cosLookup[10649] <= 0.522494477;
cosLookup[10650] <= 0.522412724;
cosLookup[10651] <= 0.522330965;
cosLookup[10652] <= 0.522249202;
cosLookup[10653] <= 0.522167434;
cosLookup[10654] <= 0.522085662;
cosLookup[10655] <= 0.522003884;
cosLookup[10656] <= 0.521922102;
cosLookup[10657] <= 0.521840315;
cosLookup[10658] <= 0.521758523;
cosLookup[10659] <= 0.521676726;
cosLookup[10660] <= 0.521594925;
cosLookup[10661] <= 0.521513119;
cosLookup[10662] <= 0.521431308;
cosLookup[10663] <= 0.521349492;
cosLookup[10664] <= 0.521267671;
cosLookup[10665] <= 0.521185846;
cosLookup[10666] <= 0.521104015;
cosLookup[10667] <= 0.52102218;
cosLookup[10668] <= 0.52094034;
cosLookup[10669] <= 0.520858496;
cosLookup[10670] <= 0.520776646;
cosLookup[10671] <= 0.520694792;
cosLookup[10672] <= 0.520612933;
cosLookup[10673] <= 0.52053107;
cosLookup[10674] <= 0.520449201;
cosLookup[10675] <= 0.520367328;
cosLookup[10676] <= 0.52028545;
cosLookup[10677] <= 0.520203567;
cosLookup[10678] <= 0.520121679;
cosLookup[10679] <= 0.520039787;
cosLookup[10680] <= 0.519957889;
cosLookup[10681] <= 0.519875987;
cosLookup[10682] <= 0.519794081;
cosLookup[10683] <= 0.519712169;
cosLookup[10684] <= 0.519630253;
cosLookup[10685] <= 0.519548332;
cosLookup[10686] <= 0.519466406;
cosLookup[10687] <= 0.519384475;
cosLookup[10688] <= 0.51930254;
cosLookup[10689] <= 0.519220599;
cosLookup[10690] <= 0.519138654;
cosLookup[10691] <= 0.519056705;
cosLookup[10692] <= 0.51897475;
cosLookup[10693] <= 0.518892791;
cosLookup[10694] <= 0.518810827;
cosLookup[10695] <= 0.518728858;
cosLookup[10696] <= 0.518646884;
cosLookup[10697] <= 0.518564906;
cosLookup[10698] <= 0.518482923;
cosLookup[10699] <= 0.518400935;
cosLookup[10700] <= 0.518318942;
cosLookup[10701] <= 0.518236945;
cosLookup[10702] <= 0.518154942;
cosLookup[10703] <= 0.518072935;
cosLookup[10704] <= 0.517990924;
cosLookup[10705] <= 0.517908907;
cosLookup[10706] <= 0.517826886;
cosLookup[10707] <= 0.51774486;
cosLookup[10708] <= 0.517662829;
cosLookup[10709] <= 0.517580794;
cosLookup[10710] <= 0.517498753;
cosLookup[10711] <= 0.517416708;
cosLookup[10712] <= 0.517334658;
cosLookup[10713] <= 0.517252604;
cosLookup[10714] <= 0.517170544;
cosLookup[10715] <= 0.51708848;
cosLookup[10716] <= 0.517006412;
cosLookup[10717] <= 0.516924338;
cosLookup[10718] <= 0.51684226;
cosLookup[10719] <= 0.516760177;
cosLookup[10720] <= 0.516678089;
cosLookup[10721] <= 0.516595996;
cosLookup[10722] <= 0.516513899;
cosLookup[10723] <= 0.516431797;
cosLookup[10724] <= 0.51634969;
cosLookup[10725] <= 0.516267578;
cosLookup[10726] <= 0.516185462;
cosLookup[10727] <= 0.516103341;
cosLookup[10728] <= 0.516021215;
cosLookup[10729] <= 0.515939084;
cosLookup[10730] <= 0.515856949;
cosLookup[10731] <= 0.515774809;
cosLookup[10732] <= 0.515692664;
cosLookup[10733] <= 0.515610515;
cosLookup[10734] <= 0.515528361;
cosLookup[10735] <= 0.515446202;
cosLookup[10736] <= 0.515364038;
cosLookup[10737] <= 0.515281869;
cosLookup[10738] <= 0.515199696;
cosLookup[10739] <= 0.515117518;
cosLookup[10740] <= 0.515035335;
cosLookup[10741] <= 0.514953148;
cosLookup[10742] <= 0.514870956;
cosLookup[10743] <= 0.514788759;
cosLookup[10744] <= 0.514706557;
cosLookup[10745] <= 0.514624351;
cosLookup[10746] <= 0.51454214;
cosLookup[10747] <= 0.514459924;
cosLookup[10748] <= 0.514377703;
cosLookup[10749] <= 0.514295478;
cosLookup[10750] <= 0.514213248;
cosLookup[10751] <= 0.514131013;
cosLookup[10752] <= 0.514048774;
cosLookup[10753] <= 0.51396653;
cosLookup[10754] <= 0.513884281;
cosLookup[10755] <= 0.513802027;
cosLookup[10756] <= 0.513719769;
cosLookup[10757] <= 0.513637506;
cosLookup[10758] <= 0.513555238;
cosLookup[10759] <= 0.513472966;
cosLookup[10760] <= 0.513390688;
cosLookup[10761] <= 0.513308406;
cosLookup[10762] <= 0.51322612;
cosLookup[10763] <= 0.513143828;
cosLookup[10764] <= 0.513061532;
cosLookup[10765] <= 0.512979231;
cosLookup[10766] <= 0.512896926;
cosLookup[10767] <= 0.512814615;
cosLookup[10768] <= 0.512732301;
cosLookup[10769] <= 0.512649981;
cosLookup[10770] <= 0.512567656;
cosLookup[10771] <= 0.512485327;
cosLookup[10772] <= 0.512402993;
cosLookup[10773] <= 0.512320655;
cosLookup[10774] <= 0.512238312;
cosLookup[10775] <= 0.512155964;
cosLookup[10776] <= 0.512073611;
cosLookup[10777] <= 0.511991254;
cosLookup[10778] <= 0.511908892;
cosLookup[10779] <= 0.511826525;
cosLookup[10780] <= 0.511744153;
cosLookup[10781] <= 0.511661777;
cosLookup[10782] <= 0.511579396;
cosLookup[10783] <= 0.511497011;
cosLookup[10784] <= 0.51141462;
cosLookup[10785] <= 0.511332225;
cosLookup[10786] <= 0.511249826;
cosLookup[10787] <= 0.511167421;
cosLookup[10788] <= 0.511085012;
cosLookup[10789] <= 0.511002598;
cosLookup[10790] <= 0.51092018;
cosLookup[10791] <= 0.510837757;
cosLookup[10792] <= 0.510755329;
cosLookup[10793] <= 0.510672896;
cosLookup[10794] <= 0.510590459;
cosLookup[10795] <= 0.510508017;
cosLookup[10796] <= 0.51042557;
cosLookup[10797] <= 0.510343119;
cosLookup[10798] <= 0.510260663;
cosLookup[10799] <= 0.510178202;
cosLookup[10800] <= 0.510095737;
cosLookup[10801] <= 0.510013267;
cosLookup[10802] <= 0.509930792;
cosLookup[10803] <= 0.509848312;
cosLookup[10804] <= 0.509765828;
cosLookup[10805] <= 0.509683339;
cosLookup[10806] <= 0.509600846;
cosLookup[10807] <= 0.509518347;
cosLookup[10808] <= 0.509435844;
cosLookup[10809] <= 0.509353337;
cosLookup[10810] <= 0.509270825;
cosLookup[10811] <= 0.509188308;
cosLookup[10812] <= 0.509105786;
cosLookup[10813] <= 0.50902326;
cosLookup[10814] <= 0.508940729;
cosLookup[10815] <= 0.508858193;
cosLookup[10816] <= 0.508775652;
cosLookup[10817] <= 0.508693107;
cosLookup[10818] <= 0.508610558;
cosLookup[10819] <= 0.508528003;
cosLookup[10820] <= 0.508445444;
cosLookup[10821] <= 0.50836288;
cosLookup[10822] <= 0.508280312;
cosLookup[10823] <= 0.508197739;
cosLookup[10824] <= 0.508115161;
cosLookup[10825] <= 0.508032579;
cosLookup[10826] <= 0.507949992;
cosLookup[10827] <= 0.5078674;
cosLookup[10828] <= 0.507784803;
cosLookup[10829] <= 0.507702202;
cosLookup[10830] <= 0.507619597;
cosLookup[10831] <= 0.507536986;
cosLookup[10832] <= 0.507454371;
cosLookup[10833] <= 0.507371751;
cosLookup[10834] <= 0.507289127;
cosLookup[10835] <= 0.507206498;
cosLookup[10836] <= 0.507123864;
cosLookup[10837] <= 0.507041225;
cosLookup[10838] <= 0.506958582;
cosLookup[10839] <= 0.506875935;
cosLookup[10840] <= 0.506793282;
cosLookup[10841] <= 0.506710625;
cosLookup[10842] <= 0.506627963;
cosLookup[10843] <= 0.506545297;
cosLookup[10844] <= 0.506462626;
cosLookup[10845] <= 0.50637995;
cosLookup[10846] <= 0.50629727;
cosLookup[10847] <= 0.506214585;
cosLookup[10848] <= 0.506131895;
cosLookup[10849] <= 0.506049201;
cosLookup[10850] <= 0.505966502;
cosLookup[10851] <= 0.505883798;
cosLookup[10852] <= 0.50580109;
cosLookup[10853] <= 0.505718377;
cosLookup[10854] <= 0.50563566;
cosLookup[10855] <= 0.505552937;
cosLookup[10856] <= 0.50547021;
cosLookup[10857] <= 0.505387479;
cosLookup[10858] <= 0.505304743;
cosLookup[10859] <= 0.505222002;
cosLookup[10860] <= 0.505139257;
cosLookup[10861] <= 0.505056506;
cosLookup[10862] <= 0.504973752;
cosLookup[10863] <= 0.504890992;
cosLookup[10864] <= 0.504808228;
cosLookup[10865] <= 0.50472546;
cosLookup[10866] <= 0.504642686;
cosLookup[10867] <= 0.504559908;
cosLookup[10868] <= 0.504477126;
cosLookup[10869] <= 0.504394339;
cosLookup[10870] <= 0.504311547;
cosLookup[10871] <= 0.50422875;
cosLookup[10872] <= 0.504145949;
cosLookup[10873] <= 0.504063143;
cosLookup[10874] <= 0.503980333;
cosLookup[10875] <= 0.503897518;
cosLookup[10876] <= 0.503814698;
cosLookup[10877] <= 0.503731874;
cosLookup[10878] <= 0.503649045;
cosLookup[10879] <= 0.503566212;
cosLookup[10880] <= 0.503483373;
cosLookup[10881] <= 0.503400531;
cosLookup[10882] <= 0.503317683;
cosLookup[10883] <= 0.503234831;
cosLookup[10884] <= 0.503151975;
cosLookup[10885] <= 0.503069113;
cosLookup[10886] <= 0.502986247;
cosLookup[10887] <= 0.502903377;
cosLookup[10888] <= 0.502820502;
cosLookup[10889] <= 0.502737622;
cosLookup[10890] <= 0.502654737;
cosLookup[10891] <= 0.502571848;
cosLookup[10892] <= 0.502488955;
cosLookup[10893] <= 0.502406056;
cosLookup[10894] <= 0.502323153;
cosLookup[10895] <= 0.502240246;
cosLookup[10896] <= 0.502157334;
cosLookup[10897] <= 0.502074417;
cosLookup[10898] <= 0.501991496;
cosLookup[10899] <= 0.50190857;
cosLookup[10900] <= 0.501825639;
cosLookup[10901] <= 0.501742704;
cosLookup[10902] <= 0.501659764;
cosLookup[10903] <= 0.50157682;
cosLookup[10904] <= 0.50149387;
cosLookup[10905] <= 0.501410917;
cosLookup[10906] <= 0.501327959;
cosLookup[10907] <= 0.501244996;
cosLookup[10908] <= 0.501162028;
cosLookup[10909] <= 0.501079056;
cosLookup[10910] <= 0.500996079;
cosLookup[10911] <= 0.500913098;
cosLookup[10912] <= 0.500830112;
cosLookup[10913] <= 0.500747122;
cosLookup[10914] <= 0.500664127;
cosLookup[10915] <= 0.500581127;
cosLookup[10916] <= 0.500498123;
cosLookup[10917] <= 0.500415114;
cosLookup[10918] <= 0.5003321;
cosLookup[10919] <= 0.500249082;
cosLookup[10920] <= 0.500166059;
cosLookup[10921] <= 0.500083032;
cosLookup[10922] <= 0.5;
cosLookup[10923] <= 0.499916963;
cosLookup[10924] <= 0.499833922;
cosLookup[10925] <= 0.499750877;
cosLookup[10926] <= 0.499667826;
cosLookup[10927] <= 0.499584771;
cosLookup[10928] <= 0.499501712;
cosLookup[10929] <= 0.499418648;
cosLookup[10930] <= 0.499335579;
cosLookup[10931] <= 0.499252506;
cosLookup[10932] <= 0.499169428;
cosLookup[10933] <= 0.499086346;
cosLookup[10934] <= 0.499003259;
cosLookup[10935] <= 0.498920167;
cosLookup[10936] <= 0.498837071;
cosLookup[10937] <= 0.49875397;
cosLookup[10938] <= 0.498670865;
cosLookup[10939] <= 0.498587755;
cosLookup[10940] <= 0.49850464;
cosLookup[10941] <= 0.498421521;
cosLookup[10942] <= 0.498338397;
cosLookup[10943] <= 0.498255269;
cosLookup[10944] <= 0.498172136;
cosLookup[10945] <= 0.498088999;
cosLookup[10946] <= 0.498005857;
cosLookup[10947] <= 0.49792271;
cosLookup[10948] <= 0.497839559;
cosLookup[10949] <= 0.497756403;
cosLookup[10950] <= 0.497673243;
cosLookup[10951] <= 0.497590078;
cosLookup[10952] <= 0.497506909;
cosLookup[10953] <= 0.497423735;
cosLookup[10954] <= 0.497340556;
cosLookup[10955] <= 0.497257373;
cosLookup[10956] <= 0.497174185;
cosLookup[10957] <= 0.497090993;
cosLookup[10958] <= 0.497007796;
cosLookup[10959] <= 0.496924594;
cosLookup[10960] <= 0.496841388;
cosLookup[10961] <= 0.496758178;
cosLookup[10962] <= 0.496674962;
cosLookup[10963] <= 0.496591743;
cosLookup[10964] <= 0.496508518;
cosLookup[10965] <= 0.49642529;
cosLookup[10966] <= 0.496342056;
cosLookup[10967] <= 0.496258818;
cosLookup[10968] <= 0.496175576;
cosLookup[10969] <= 0.496092328;
cosLookup[10970] <= 0.496009077;
cosLookup[10971] <= 0.49592582;
cosLookup[10972] <= 0.49584256;
cosLookup[10973] <= 0.495759294;
cosLookup[10974] <= 0.495676024;
cosLookup[10975] <= 0.49559275;
cosLookup[10976] <= 0.495509471;
cosLookup[10977] <= 0.495426187;
cosLookup[10978] <= 0.495342899;
cosLookup[10979] <= 0.495259606;
cosLookup[10980] <= 0.495176309;
cosLookup[10981] <= 0.495093007;
cosLookup[10982] <= 0.495009701;
cosLookup[10983] <= 0.49492639;
cosLookup[10984] <= 0.494843075;
cosLookup[10985] <= 0.494759755;
cosLookup[10986] <= 0.49467643;
cosLookup[10987] <= 0.494593101;
cosLookup[10988] <= 0.494509767;
cosLookup[10989] <= 0.494426429;
cosLookup[10990] <= 0.494343087;
cosLookup[10991] <= 0.494259739;
cosLookup[10992] <= 0.494176387;
cosLookup[10993] <= 0.494093031;
cosLookup[10994] <= 0.49400967;
cosLookup[10995] <= 0.493926305;
cosLookup[10996] <= 0.493842935;
cosLookup[10997] <= 0.49375956;
cosLookup[10998] <= 0.493676181;
cosLookup[10999] <= 0.493592797;
cosLookup[11000] <= 0.493509409;
cosLookup[11001] <= 0.493426017;
cosLookup[11002] <= 0.493342619;
cosLookup[11003] <= 0.493259218;
cosLookup[11004] <= 0.493175811;
cosLookup[11005] <= 0.493092401;
cosLookup[11006] <= 0.493008985;
cosLookup[11007] <= 0.492925565;
cosLookup[11008] <= 0.492842141;
cosLookup[11009] <= 0.492758712;
cosLookup[11010] <= 0.492675279;
cosLookup[11011] <= 0.492591841;
cosLookup[11012] <= 0.492508398;
cosLookup[11013] <= 0.492424951;
cosLookup[11014] <= 0.492341499;
cosLookup[11015] <= 0.492258043;
cosLookup[11016] <= 0.492174583;
cosLookup[11017] <= 0.492091117;
cosLookup[11018] <= 0.492007648;
cosLookup[11019] <= 0.491924174;
cosLookup[11020] <= 0.491840695;
cosLookup[11021] <= 0.491757212;
cosLookup[11022] <= 0.491673724;
cosLookup[11023] <= 0.491590231;
cosLookup[11024] <= 0.491506735;
cosLookup[11025] <= 0.491423233;
cosLookup[11026] <= 0.491339727;
cosLookup[11027] <= 0.491256217;
cosLookup[11028] <= 0.491172702;
cosLookup[11029] <= 0.491089183;
cosLookup[11030] <= 0.491005659;
cosLookup[11031] <= 0.49092213;
cosLookup[11032] <= 0.490838598;
cosLookup[11033] <= 0.49075506;
cosLookup[11034] <= 0.490671518;
cosLookup[11035] <= 0.490587972;
cosLookup[11036] <= 0.490504421;
cosLookup[11037] <= 0.490420865;
cosLookup[11038] <= 0.490337305;
cosLookup[11039] <= 0.490253741;
cosLookup[11040] <= 0.490170172;
cosLookup[11041] <= 0.490086598;
cosLookup[11042] <= 0.49000302;
cosLookup[11043] <= 0.489919438;
cosLookup[11044] <= 0.489835851;
cosLookup[11045] <= 0.489752259;
cosLookup[11046] <= 0.489668663;
cosLookup[11047] <= 0.489585062;
cosLookup[11048] <= 0.489501457;
cosLookup[11049] <= 0.489417848;
cosLookup[11050] <= 0.489334234;
cosLookup[11051] <= 0.489250615;
cosLookup[11052] <= 0.489166992;
cosLookup[11053] <= 0.489083365;
cosLookup[11054] <= 0.488999733;
cosLookup[11055] <= 0.488916096;
cosLookup[11056] <= 0.488832455;
cosLookup[11057] <= 0.48874881;
cosLookup[11058] <= 0.48866516;
cosLookup[11059] <= 0.488581505;
cosLookup[11060] <= 0.488497846;
cosLookup[11061] <= 0.488414183;
cosLookup[11062] <= 0.488330515;
cosLookup[11063] <= 0.488246842;
cosLookup[11064] <= 0.488163165;
cosLookup[11065] <= 0.488079484;
cosLookup[11066] <= 0.487995798;
cosLookup[11067] <= 0.487912107;
cosLookup[11068] <= 0.487828413;
cosLookup[11069] <= 0.487744713;
cosLookup[11070] <= 0.487661009;
cosLookup[11071] <= 0.487577301;
cosLookup[11072] <= 0.487493588;
cosLookup[11073] <= 0.487409871;
cosLookup[11074] <= 0.487326149;
cosLookup[11075] <= 0.487242423;
cosLookup[11076] <= 0.487158692;
cosLookup[11077] <= 0.487074957;
cosLookup[11078] <= 0.486991217;
cosLookup[11079] <= 0.486907473;
cosLookup[11080] <= 0.486823724;
cosLookup[11081] <= 0.486739971;
cosLookup[11082] <= 0.486656213;
cosLookup[11083] <= 0.486572451;
cosLookup[11084] <= 0.486488685;
cosLookup[11085] <= 0.486404914;
cosLookup[11086] <= 0.486321138;
cosLookup[11087] <= 0.486237358;
cosLookup[11088] <= 0.486153574;
cosLookup[11089] <= 0.486069785;
cosLookup[11090] <= 0.485985992;
cosLookup[11091] <= 0.485902194;
cosLookup[11092] <= 0.485818391;
cosLookup[11093] <= 0.485734585;
cosLookup[11094] <= 0.485650773;
cosLookup[11095] <= 0.485566958;
cosLookup[11096] <= 0.485483138;
cosLookup[11097] <= 0.485399313;
cosLookup[11098] <= 0.485315484;
cosLookup[11099] <= 0.48523165;
cosLookup[11100] <= 0.485147812;
cosLookup[11101] <= 0.48506397;
cosLookup[11102] <= 0.484980123;
cosLookup[11103] <= 0.484896271;
cosLookup[11104] <= 0.484812416;
cosLookup[11105] <= 0.484728555;
cosLookup[11106] <= 0.48464469;
cosLookup[11107] <= 0.484560821;
cosLookup[11108] <= 0.484476948;
cosLookup[11109] <= 0.484393069;
cosLookup[11110] <= 0.484309187;
cosLookup[11111] <= 0.4842253;
cosLookup[11112] <= 0.484141408;
cosLookup[11113] <= 0.484057512;
cosLookup[11114] <= 0.483973612;
cosLookup[11115] <= 0.483889707;
cosLookup[11116] <= 0.483805798;
cosLookup[11117] <= 0.483721884;
cosLookup[11118] <= 0.483637966;
cosLookup[11119] <= 0.483554043;
cosLookup[11120] <= 0.483470116;
cosLookup[11121] <= 0.483386185;
cosLookup[11122] <= 0.483302249;
cosLookup[11123] <= 0.483218308;
cosLookup[11124] <= 0.483134364;
cosLookup[11125] <= 0.483050414;
cosLookup[11126] <= 0.48296646;
cosLookup[11127] <= 0.482882502;
cosLookup[11128] <= 0.48279854;
cosLookup[11129] <= 0.482714573;
cosLookup[11130] <= 0.482630601;
cosLookup[11131] <= 0.482546625;
cosLookup[11132] <= 0.482462645;
cosLookup[11133] <= 0.48237866;
cosLookup[11134] <= 0.482294671;
cosLookup[11135] <= 0.482210677;
cosLookup[11136] <= 0.482126679;
cosLookup[11137] <= 0.482042677;
cosLookup[11138] <= 0.48195867;
cosLookup[11139] <= 0.481874658;
cosLookup[11140] <= 0.481790642;
cosLookup[11141] <= 0.481706622;
cosLookup[11142] <= 0.481622598;
cosLookup[11143] <= 0.481538568;
cosLookup[11144] <= 0.481454535;
cosLookup[11145] <= 0.481370497;
cosLookup[11146] <= 0.481286455;
cosLookup[11147] <= 0.481202408;
cosLookup[11148] <= 0.481118357;
cosLookup[11149] <= 0.481034301;
cosLookup[11150] <= 0.480950241;
cosLookup[11151] <= 0.480866176;
cosLookup[11152] <= 0.480782107;
cosLookup[11153] <= 0.480698034;
cosLookup[11154] <= 0.480613956;
cosLookup[11155] <= 0.480529874;
cosLookup[11156] <= 0.480445788;
cosLookup[11157] <= 0.480361697;
cosLookup[11158] <= 0.480277601;
cosLookup[11159] <= 0.480193501;
cosLookup[11160] <= 0.480109397;
cosLookup[11161] <= 0.480025288;
cosLookup[11162] <= 0.479941175;
cosLookup[11163] <= 0.479857058;
cosLookup[11164] <= 0.479772936;
cosLookup[11165] <= 0.47968881;
cosLookup[11166] <= 0.479604679;
cosLookup[11167] <= 0.479520544;
cosLookup[11168] <= 0.479436404;
cosLookup[11169] <= 0.47935226;
cosLookup[11170] <= 0.479268112;
cosLookup[11171] <= 0.479183959;
cosLookup[11172] <= 0.479099802;
cosLookup[11173] <= 0.47901564;
cosLookup[11174] <= 0.478931475;
cosLookup[11175] <= 0.478847304;
cosLookup[11176] <= 0.478763129;
cosLookup[11177] <= 0.47867895;
cosLookup[11178] <= 0.478594767;
cosLookup[11179] <= 0.478510579;
cosLookup[11180] <= 0.478426386;
cosLookup[11181] <= 0.478342189;
cosLookup[11182] <= 0.478257988;
cosLookup[11183] <= 0.478173783;
cosLookup[11184] <= 0.478089573;
cosLookup[11185] <= 0.478005358;
cosLookup[11186] <= 0.47792114;
cosLookup[11187] <= 0.477836917;
cosLookup[11188] <= 0.477752689;
cosLookup[11189] <= 0.477668457;
cosLookup[11190] <= 0.477584221;
cosLookup[11191] <= 0.47749998;
cosLookup[11192] <= 0.477415735;
cosLookup[11193] <= 0.477331485;
cosLookup[11194] <= 0.477247232;
cosLookup[11195] <= 0.477162973;
cosLookup[11196] <= 0.477078711;
cosLookup[11197] <= 0.476994444;
cosLookup[11198] <= 0.476910172;
cosLookup[11199] <= 0.476825896;
cosLookup[11200] <= 0.476741616;
cosLookup[11201] <= 0.476657332;
cosLookup[11202] <= 0.476573043;
cosLookup[11203] <= 0.476488749;
cosLookup[11204] <= 0.476404452;
cosLookup[11205] <= 0.47632015;
cosLookup[11206] <= 0.476235843;
cosLookup[11207] <= 0.476151532;
cosLookup[11208] <= 0.476067217;
cosLookup[11209] <= 0.475982897;
cosLookup[11210] <= 0.475898573;
cosLookup[11211] <= 0.475814245;
cosLookup[11212] <= 0.475729912;
cosLookup[11213] <= 0.475645575;
cosLookup[11214] <= 0.475561234;
cosLookup[11215] <= 0.475476888;
cosLookup[11216] <= 0.475392538;
cosLookup[11217] <= 0.475308183;
cosLookup[11218] <= 0.475223824;
cosLookup[11219] <= 0.475139461;
cosLookup[11220] <= 0.475055093;
cosLookup[11221] <= 0.474970721;
cosLookup[11222] <= 0.474886345;
cosLookup[11223] <= 0.474801964;
cosLookup[11224] <= 0.474717579;
cosLookup[11225] <= 0.474633189;
cosLookup[11226] <= 0.474548795;
cosLookup[11227] <= 0.474464397;
cosLookup[11228] <= 0.474379994;
cosLookup[11229] <= 0.474295587;
cosLookup[11230] <= 0.474211176;
cosLookup[11231] <= 0.47412676;
cosLookup[11232] <= 0.47404234;
cosLookup[11233] <= 0.473957916;
cosLookup[11234] <= 0.473873487;
cosLookup[11235] <= 0.473789054;
cosLookup[11236] <= 0.473704617;
cosLookup[11237] <= 0.473620175;
cosLookup[11238] <= 0.473535728;
cosLookup[11239] <= 0.473451278;
cosLookup[11240] <= 0.473366823;
cosLookup[11241] <= 0.473282364;
cosLookup[11242] <= 0.4731979;
cosLookup[11243] <= 0.473113432;
cosLookup[11244] <= 0.47302896;
cosLookup[11245] <= 0.472944483;
cosLookup[11246] <= 0.472860002;
cosLookup[11247] <= 0.472775517;
cosLookup[11248] <= 0.472691027;
cosLookup[11249] <= 0.472606533;
cosLookup[11250] <= 0.472522035;
cosLookup[11251] <= 0.472437532;
cosLookup[11252] <= 0.472353025;
cosLookup[11253] <= 0.472268514;
cosLookup[11254] <= 0.472183998;
cosLookup[11255] <= 0.472099478;
cosLookup[11256] <= 0.472014954;
cosLookup[11257] <= 0.471930425;
cosLookup[11258] <= 0.471845892;
cosLookup[11259] <= 0.471761354;
cosLookup[11260] <= 0.471676812;
cosLookup[11261] <= 0.471592266;
cosLookup[11262] <= 0.471507716;
cosLookup[11263] <= 0.471423161;
cosLookup[11264] <= 0.471338602;
cosLookup[11265] <= 0.471254039;
cosLookup[11266] <= 0.471169471;
cosLookup[11267] <= 0.471084899;
cosLookup[11268] <= 0.471000322;
cosLookup[11269] <= 0.470915741;
cosLookup[11270] <= 0.470831156;
cosLookup[11271] <= 0.470746567;
cosLookup[11272] <= 0.470661973;
cosLookup[11273] <= 0.470577375;
cosLookup[11274] <= 0.470492773;
cosLookup[11275] <= 0.470408166;
cosLookup[11276] <= 0.470323555;
cosLookup[11277] <= 0.470238939;
cosLookup[11278] <= 0.47015432;
cosLookup[11279] <= 0.470069696;
cosLookup[11280] <= 0.469985067;
cosLookup[11281] <= 0.469900435;
cosLookup[11282] <= 0.469815798;
cosLookup[11283] <= 0.469731156;
cosLookup[11284] <= 0.469646511;
cosLookup[11285] <= 0.469561861;
cosLookup[11286] <= 0.469477207;
cosLookup[11287] <= 0.469392548;
cosLookup[11288] <= 0.469307885;
cosLookup[11289] <= 0.469223218;
cosLookup[11290] <= 0.469138546;
cosLookup[11291] <= 0.469053871;
cosLookup[11292] <= 0.46896919;
cosLookup[11293] <= 0.468884506;
cosLookup[11294] <= 0.468799817;
cosLookup[11295] <= 0.468715124;
cosLookup[11296] <= 0.468630427;
cosLookup[11297] <= 0.468545725;
cosLookup[11298] <= 0.468461019;
cosLookup[11299] <= 0.468376309;
cosLookup[11300] <= 0.468291594;
cosLookup[11301] <= 0.468206875;
cosLookup[11302] <= 0.468122152;
cosLookup[11303] <= 0.468037424;
cosLookup[11304] <= 0.467952693;
cosLookup[11305] <= 0.467867956;
cosLookup[11306] <= 0.467783216;
cosLookup[11307] <= 0.467698471;
cosLookup[11308] <= 0.467613722;
cosLookup[11309] <= 0.467528969;
cosLookup[11310] <= 0.467444211;
cosLookup[11311] <= 0.467359449;
cosLookup[11312] <= 0.467274683;
cosLookup[11313] <= 0.467189913;
cosLookup[11314] <= 0.467105138;
cosLookup[11315] <= 0.467020359;
cosLookup[11316] <= 0.466935575;
cosLookup[11317] <= 0.466850788;
cosLookup[11318] <= 0.466765996;
cosLookup[11319] <= 0.466681199;
cosLookup[11320] <= 0.466596399;
cosLookup[11321] <= 0.466511594;
cosLookup[11322] <= 0.466426785;
cosLookup[11323] <= 0.466341971;
cosLookup[11324] <= 0.466257154;
cosLookup[11325] <= 0.466172332;
cosLookup[11326] <= 0.466087505;
cosLookup[11327] <= 0.466002675;
cosLookup[11328] <= 0.46591784;
cosLookup[11329] <= 0.465833001;
cosLookup[11330] <= 0.465748157;
cosLookup[11331] <= 0.46566331;
cosLookup[11332] <= 0.465578458;
cosLookup[11333] <= 0.465493601;
cosLookup[11334] <= 0.465408741;
cosLookup[11335] <= 0.465323876;
cosLookup[11336] <= 0.465239007;
cosLookup[11337] <= 0.465154134;
cosLookup[11338] <= 0.465069256;
cosLookup[11339] <= 0.464984374;
cosLookup[11340] <= 0.464899488;
cosLookup[11341] <= 0.464814597;
cosLookup[11342] <= 0.464729703;
cosLookup[11343] <= 0.464644804;
cosLookup[11344] <= 0.4645599;
cosLookup[11345] <= 0.464474993;
cosLookup[11346] <= 0.464390081;
cosLookup[11347] <= 0.464305165;
cosLookup[11348] <= 0.464220244;
cosLookup[11349] <= 0.46413532;
cosLookup[11350] <= 0.464050391;
cosLookup[11351] <= 0.463965458;
cosLookup[11352] <= 0.46388052;
cosLookup[11353] <= 0.463795579;
cosLookup[11354] <= 0.463710633;
cosLookup[11355] <= 0.463625682;
cosLookup[11356] <= 0.463540728;
cosLookup[11357] <= 0.463455769;
cosLookup[11358] <= 0.463370806;
cosLookup[11359] <= 0.463285839;
cosLookup[11360] <= 0.463200867;
cosLookup[11361] <= 0.463115892;
cosLookup[11362] <= 0.463030911;
cosLookup[11363] <= 0.462945927;
cosLookup[11364] <= 0.462860939;
cosLookup[11365] <= 0.462775946;
cosLookup[11366] <= 0.462690949;
cosLookup[11367] <= 0.462605947;
cosLookup[11368] <= 0.462520942;
cosLookup[11369] <= 0.462435932;
cosLookup[11370] <= 0.462350918;
cosLookup[11371] <= 0.4622659;
cosLookup[11372] <= 0.462180877;
cosLookup[11373] <= 0.46209585;
cosLookup[11374] <= 0.462010819;
cosLookup[11375] <= 0.461925784;
cosLookup[11376] <= 0.461840744;
cosLookup[11377] <= 0.4617557;
cosLookup[11378] <= 0.461670652;
cosLookup[11379] <= 0.4615856;
cosLookup[11380] <= 0.461500544;
cosLookup[11381] <= 0.461415483;
cosLookup[11382] <= 0.461330418;
cosLookup[11383] <= 0.461245348;
cosLookup[11384] <= 0.461160275;
cosLookup[11385] <= 0.461075197;
cosLookup[11386] <= 0.460990115;
cosLookup[11387] <= 0.460905029;
cosLookup[11388] <= 0.460819938;
cosLookup[11389] <= 0.460734844;
cosLookup[11390] <= 0.460649745;
cosLookup[11391] <= 0.460564642;
cosLookup[11392] <= 0.460479534;
cosLookup[11393] <= 0.460394423;
cosLookup[11394] <= 0.460309307;
cosLookup[11395] <= 0.460224187;
cosLookup[11396] <= 0.460139062;
cosLookup[11397] <= 0.460053934;
cosLookup[11398] <= 0.459968801;
cosLookup[11399] <= 0.459883664;
cosLookup[11400] <= 0.459798523;
cosLookup[11401] <= 0.459713377;
cosLookup[11402] <= 0.459628228;
cosLookup[11403] <= 0.459543074;
cosLookup[11404] <= 0.459457915;
cosLookup[11405] <= 0.459372753;
cosLookup[11406] <= 0.459287586;
cosLookup[11407] <= 0.459202416;
cosLookup[11408] <= 0.459117241;
cosLookup[11409] <= 0.459032061;
cosLookup[11410] <= 0.458946878;
cosLookup[11411] <= 0.45886169;
cosLookup[11412] <= 0.458776498;
cosLookup[11413] <= 0.458691302;
cosLookup[11414] <= 0.458606102;
cosLookup[11415] <= 0.458520897;
cosLookup[11416] <= 0.458435688;
cosLookup[11417] <= 0.458350475;
cosLookup[11418] <= 0.458265258;
cosLookup[11419] <= 0.458180037;
cosLookup[11420] <= 0.458094811;
cosLookup[11421] <= 0.458009581;
cosLookup[11422] <= 0.457924347;
cosLookup[11423] <= 0.457839109;
cosLookup[11424] <= 0.457753867;
cosLookup[11425] <= 0.45766862;
cosLookup[11426] <= 0.457583369;
cosLookup[11427] <= 0.457498114;
cosLookup[11428] <= 0.457412855;
cosLookup[11429] <= 0.457327591;
cosLookup[11430] <= 0.457242323;
cosLookup[11431] <= 0.457157051;
cosLookup[11432] <= 0.457071775;
cosLookup[11433] <= 0.456986495;
cosLookup[11434] <= 0.45690121;
cosLookup[11435] <= 0.456815922;
cosLookup[11436] <= 0.456730629;
cosLookup[11437] <= 0.456645332;
cosLookup[11438] <= 0.45656003;
cosLookup[11439] <= 0.456474725;
cosLookup[11440] <= 0.456389415;
cosLookup[11441] <= 0.456304101;
cosLookup[11442] <= 0.456218783;
cosLookup[11443] <= 0.456133461;
cosLookup[11444] <= 0.456048134;
cosLookup[11445] <= 0.455962804;
cosLookup[11446] <= 0.455877469;
cosLookup[11447] <= 0.45579213;
cosLookup[11448] <= 0.455706786;
cosLookup[11449] <= 0.455621439;
cosLookup[11450] <= 0.455536087;
cosLookup[11451] <= 0.455450732;
cosLookup[11452] <= 0.455365372;
cosLookup[11453] <= 0.455280007;
cosLookup[11454] <= 0.455194639;
cosLookup[11455] <= 0.455109266;
cosLookup[11456] <= 0.45502389;
cosLookup[11457] <= 0.454938509;
cosLookup[11458] <= 0.454853124;
cosLookup[11459] <= 0.454767734;
cosLookup[11460] <= 0.454682341;
cosLookup[11461] <= 0.454596943;
cosLookup[11462] <= 0.454511541;
cosLookup[11463] <= 0.454426135;
cosLookup[11464] <= 0.454340725;
cosLookup[11465] <= 0.454255311;
cosLookup[11466] <= 0.454169892;
cosLookup[11467] <= 0.45408447;
cosLookup[11468] <= 0.453999043;
cosLookup[11469] <= 0.453913612;
cosLookup[11470] <= 0.453828176;
cosLookup[11471] <= 0.453742737;
cosLookup[11472] <= 0.453657293;
cosLookup[11473] <= 0.453571846;
cosLookup[11474] <= 0.453486394;
cosLookup[11475] <= 0.453400938;
cosLookup[11476] <= 0.453315477;
cosLookup[11477] <= 0.453230013;
cosLookup[11478] <= 0.453144544;
cosLookup[11479] <= 0.453059072;
cosLookup[11480] <= 0.452973595;
cosLookup[11481] <= 0.452888114;
cosLookup[11482] <= 0.452802628;
cosLookup[11483] <= 0.452717139;
cosLookup[11484] <= 0.452631645;
cosLookup[11485] <= 0.452546148;
cosLookup[11486] <= 0.452460646;
cosLookup[11487] <= 0.45237514;
cosLookup[11488] <= 0.452289629;
cosLookup[11489] <= 0.452204115;
cosLookup[11490] <= 0.452118597;
cosLookup[11491] <= 0.452033074;
cosLookup[11492] <= 0.451947547;
cosLookup[11493] <= 0.451862016;
cosLookup[11494] <= 0.451776481;
cosLookup[11495] <= 0.451690942;
cosLookup[11496] <= 0.451605398;
cosLookup[11497] <= 0.451519851;
cosLookup[11498] <= 0.451434299;
cosLookup[11499] <= 0.451348743;
cosLookup[11500] <= 0.451263183;
cosLookup[11501] <= 0.451177619;
cosLookup[11502] <= 0.45109205;
cosLookup[11503] <= 0.451006478;
cosLookup[11504] <= 0.450920901;
cosLookup[11505] <= 0.45083532;
cosLookup[11506] <= 0.450749735;
cosLookup[11507] <= 0.450664146;
cosLookup[11508] <= 0.450578553;
cosLookup[11509] <= 0.450492956;
cosLookup[11510] <= 0.450407354;
cosLookup[11511] <= 0.450321749;
cosLookup[11512] <= 0.450236139;
cosLookup[11513] <= 0.450150525;
cosLookup[11514] <= 0.450064907;
cosLookup[11515] <= 0.449979285;
cosLookup[11516] <= 0.449893658;
cosLookup[11517] <= 0.449808028;
cosLookup[11518] <= 0.449722393;
cosLookup[11519] <= 0.449636754;
cosLookup[11520] <= 0.449551112;
cosLookup[11521] <= 0.449465465;
cosLookup[11522] <= 0.449379813;
cosLookup[11523] <= 0.449294158;
cosLookup[11524] <= 0.449208499;
cosLookup[11525] <= 0.449122835;
cosLookup[11526] <= 0.449037168;
cosLookup[11527] <= 0.448951496;
cosLookup[11528] <= 0.44886582;
cosLookup[11529] <= 0.44878014;
cosLookup[11530] <= 0.448694456;
cosLookup[11531] <= 0.448608767;
cosLookup[11532] <= 0.448523075;
cosLookup[11533] <= 0.448437378;
cosLookup[11534] <= 0.448351678;
cosLookup[11535] <= 0.448265973;
cosLookup[11536] <= 0.448180264;
cosLookup[11537] <= 0.448094551;
cosLookup[11538] <= 0.448008834;
cosLookup[11539] <= 0.447923113;
cosLookup[11540] <= 0.447837387;
cosLookup[11541] <= 0.447751658;
cosLookup[11542] <= 0.447665924;
cosLookup[11543] <= 0.447580186;
cosLookup[11544] <= 0.447494445;
cosLookup[11545] <= 0.447408699;
cosLookup[11546] <= 0.447322949;
cosLookup[11547] <= 0.447237194;
cosLookup[11548] <= 0.447151436;
cosLookup[11549] <= 0.447065674;
cosLookup[11550] <= 0.446979907;
cosLookup[11551] <= 0.446894137;
cosLookup[11552] <= 0.446808362;
cosLookup[11553] <= 0.446722583;
cosLookup[11554] <= 0.4466368;
cosLookup[11555] <= 0.446551013;
cosLookup[11556] <= 0.446465222;
cosLookup[11557] <= 0.446379427;
cosLookup[11558] <= 0.446293627;
cosLookup[11559] <= 0.446207824;
cosLookup[11560] <= 0.446122016;
cosLookup[11561] <= 0.446036205;
cosLookup[11562] <= 0.445950389;
cosLookup[11563] <= 0.445864569;
cosLookup[11564] <= 0.445778745;
cosLookup[11565] <= 0.445692917;
cosLookup[11566] <= 0.445607085;
cosLookup[11567] <= 0.445521248;
cosLookup[11568] <= 0.445435408;
cosLookup[11569] <= 0.445349564;
cosLookup[11570] <= 0.445263715;
cosLookup[11571] <= 0.445177862;
cosLookup[11572] <= 0.445092006;
cosLookup[11573] <= 0.445006145;
cosLookup[11574] <= 0.44492028;
cosLookup[11575] <= 0.444834411;
cosLookup[11576] <= 0.444748538;
cosLookup[11577] <= 0.444662661;
cosLookup[11578] <= 0.444576779;
cosLookup[11579] <= 0.444490894;
cosLookup[11580] <= 0.444405005;
cosLookup[11581] <= 0.444319111;
cosLookup[11582] <= 0.444233214;
cosLookup[11583] <= 0.444147312;
cosLookup[11584] <= 0.444061406;
cosLookup[11585] <= 0.443975496;
cosLookup[11586] <= 0.443889582;
cosLookup[11587] <= 0.443803664;
cosLookup[11588] <= 0.443717742;
cosLookup[11589] <= 0.443631816;
cosLookup[11590] <= 0.443545886;
cosLookup[11591] <= 0.443459951;
cosLookup[11592] <= 0.443374013;
cosLookup[11593] <= 0.44328807;
cosLookup[11594] <= 0.443202124;
cosLookup[11595] <= 0.443116173;
cosLookup[11596] <= 0.443030219;
cosLookup[11597] <= 0.44294426;
cosLookup[11598] <= 0.442858297;
cosLookup[11599] <= 0.44277233;
cosLookup[11600] <= 0.442686359;
cosLookup[11601] <= 0.442600384;
cosLookup[11602] <= 0.442514405;
cosLookup[11603] <= 0.442428422;
cosLookup[11604] <= 0.442342434;
cosLookup[11605] <= 0.442256443;
cosLookup[11606] <= 0.442170448;
cosLookup[11607] <= 0.442084448;
cosLookup[11608] <= 0.441998445;
cosLookup[11609] <= 0.441912437;
cosLookup[11610] <= 0.441826425;
cosLookup[11611] <= 0.44174041;
cosLookup[11612] <= 0.44165439;
cosLookup[11613] <= 0.441568366;
cosLookup[11614] <= 0.441482338;
cosLookup[11615] <= 0.441396306;
cosLookup[11616] <= 0.44131027;
cosLookup[11617] <= 0.44122423;
cosLookup[11618] <= 0.441138186;
cosLookup[11619] <= 0.441052138;
cosLookup[11620] <= 0.440966085;
cosLookup[11621] <= 0.440880029;
cosLookup[11622] <= 0.440793969;
cosLookup[11623] <= 0.440707904;
cosLookup[11624] <= 0.440621836;
cosLookup[11625] <= 0.440535764;
cosLookup[11626] <= 0.440449687;
cosLookup[11627] <= 0.440363606;
cosLookup[11628] <= 0.440277522;
cosLookup[11629] <= 0.440191433;
cosLookup[11630] <= 0.44010534;
cosLookup[11631] <= 0.440019243;
cosLookup[11632] <= 0.439933143;
cosLookup[11633] <= 0.439847038;
cosLookup[11634] <= 0.439760929;
cosLookup[11635] <= 0.439674816;
cosLookup[11636] <= 0.439588699;
cosLookup[11637] <= 0.439502578;
cosLookup[11638] <= 0.439416453;
cosLookup[11639] <= 0.439330324;
cosLookup[11640] <= 0.43924419;
cosLookup[11641] <= 0.439158053;
cosLookup[11642] <= 0.439071912;
cosLookup[11643] <= 0.438985767;
cosLookup[11644] <= 0.438899617;
cosLookup[11645] <= 0.438813464;
cosLookup[11646] <= 0.438727307;
cosLookup[11647] <= 0.438641145;
cosLookup[11648] <= 0.43855498;
cosLookup[11649] <= 0.43846881;
cosLookup[11650] <= 0.438382637;
cosLookup[11651] <= 0.438296459;
cosLookup[11652] <= 0.438210278;
cosLookup[11653] <= 0.438124092;
cosLookup[11654] <= 0.438037903;
cosLookup[11655] <= 0.437951709;
cosLookup[11656] <= 0.437865511;
cosLookup[11657] <= 0.43777931;
cosLookup[11658] <= 0.437693104;
cosLookup[11659] <= 0.437606894;
cosLookup[11660] <= 0.43752068;
cosLookup[11661] <= 0.437434463;
cosLookup[11662] <= 0.437348241;
cosLookup[11663] <= 0.437262015;
cosLookup[11664] <= 0.437175785;
cosLookup[11665] <= 0.437089551;
cosLookup[11666] <= 0.437003313;
cosLookup[11667] <= 0.436917071;
cosLookup[11668] <= 0.436830825;
cosLookup[11669] <= 0.436744575;
cosLookup[11670] <= 0.436658322;
cosLookup[11671] <= 0.436572064;
cosLookup[11672] <= 0.436485802;
cosLookup[11673] <= 0.436399536;
cosLookup[11674] <= 0.436313266;
cosLookup[11675] <= 0.436226992;
cosLookup[11676] <= 0.436140713;
cosLookup[11677] <= 0.436054431;
cosLookup[11678] <= 0.435968145;
cosLookup[11679] <= 0.435881855;
cosLookup[11680] <= 0.435795561;
cosLookup[11681] <= 0.435709263;
cosLookup[11682] <= 0.435622961;
cosLookup[11683] <= 0.435536655;
cosLookup[11684] <= 0.435450345;
cosLookup[11685] <= 0.435364031;
cosLookup[11686] <= 0.435277713;
cosLookup[11687] <= 0.435191391;
cosLookup[11688] <= 0.435105065;
cosLookup[11689] <= 0.435018735;
cosLookup[11690] <= 0.4349324;
cosLookup[11691] <= 0.434846062;
cosLookup[11692] <= 0.43475972;
cosLookup[11693] <= 0.434673374;
cosLookup[11694] <= 0.434587024;
cosLookup[11695] <= 0.43450067;
cosLookup[11696] <= 0.434414312;
cosLookup[11697] <= 0.43432795;
cosLookup[11698] <= 0.434241584;
cosLookup[11699] <= 0.434155214;
cosLookup[11700] <= 0.43406884;
cosLookup[11701] <= 0.433982462;
cosLookup[11702] <= 0.43389608;
cosLookup[11703] <= 0.433809694;
cosLookup[11704] <= 0.433723304;
cosLookup[11705] <= 0.43363691;
cosLookup[11706] <= 0.433550512;
cosLookup[11707] <= 0.43346411;
cosLookup[11708] <= 0.433377704;
cosLookup[11709] <= 0.433291294;
cosLookup[11710] <= 0.43320488;
cosLookup[11711] <= 0.433118462;
cosLookup[11712] <= 0.43303204;
cosLookup[11713] <= 0.432945614;
cosLookup[11714] <= 0.432859185;
cosLookup[11715] <= 0.432772751;
cosLookup[11716] <= 0.432686313;
cosLookup[11717] <= 0.432599871;
cosLookup[11718] <= 0.432513426;
cosLookup[11719] <= 0.432426976;
cosLookup[11720] <= 0.432340522;
cosLookup[11721] <= 0.432254064;
cosLookup[11722] <= 0.432167603;
cosLookup[11723] <= 0.432081137;
cosLookup[11724] <= 0.431994668;
cosLookup[11725] <= 0.431908194;
cosLookup[11726] <= 0.431821717;
cosLookup[11727] <= 0.431735235;
cosLookup[11728] <= 0.43164875;
cosLookup[11729] <= 0.43156226;
cosLookup[11730] <= 0.431475767;
cosLookup[11731] <= 0.431389269;
cosLookup[11732] <= 0.431302768;
cosLookup[11733] <= 0.431216263;
cosLookup[11734] <= 0.431129753;
cosLookup[11735] <= 0.43104324;
cosLookup[11736] <= 0.430956723;
cosLookup[11737] <= 0.430870202;
cosLookup[11738] <= 0.430783677;
cosLookup[11739] <= 0.430697148;
cosLookup[11740] <= 0.430610615;
cosLookup[11741] <= 0.430524078;
cosLookup[11742] <= 0.430437537;
cosLookup[11743] <= 0.430350992;
cosLookup[11744] <= 0.430264443;
cosLookup[11745] <= 0.43017789;
cosLookup[11746] <= 0.430091333;
cosLookup[11747] <= 0.430004773;
cosLookup[11748] <= 0.429918208;
cosLookup[11749] <= 0.429831639;
cosLookup[11750] <= 0.429745067;
cosLookup[11751] <= 0.42965849;
cosLookup[11752] <= 0.42957191;
cosLookup[11753] <= 0.429485325;
cosLookup[11754] <= 0.429398737;
cosLookup[11755] <= 0.429312145;
cosLookup[11756] <= 0.429225548;
cosLookup[11757] <= 0.429138948;
cosLookup[11758] <= 0.429052344;
cosLookup[11759] <= 0.428965736;
cosLookup[11760] <= 0.428879124;
cosLookup[11761] <= 0.428792508;
cosLookup[11762] <= 0.428705888;
cosLookup[11763] <= 0.428619264;
cosLookup[11764] <= 0.428532636;
cosLookup[11765] <= 0.428446004;
cosLookup[11766] <= 0.428359369;
cosLookup[11767] <= 0.428272729;
cosLookup[11768] <= 0.428186086;
cosLookup[11769] <= 0.428099438;
cosLookup[11770] <= 0.428012787;
cosLookup[11771] <= 0.427926131;
cosLookup[11772] <= 0.427839472;
cosLookup[11773] <= 0.427752809;
cosLookup[11774] <= 0.427666141;
cosLookup[11775] <= 0.42757947;
cosLookup[11776] <= 0.427492795;
cosLookup[11777] <= 0.427406116;
cosLookup[11778] <= 0.427319433;
cosLookup[11779] <= 0.427232747;
cosLookup[11780] <= 0.427146056;
cosLookup[11781] <= 0.427059361;
cosLookup[11782] <= 0.426972663;
cosLookup[11783] <= 0.42688596;
cosLookup[11784] <= 0.426799254;
cosLookup[11785] <= 0.426712543;
cosLookup[11786] <= 0.426625829;
cosLookup[11787] <= 0.426539111;
cosLookup[11788] <= 0.426452389;
cosLookup[11789] <= 0.426365663;
cosLookup[11790] <= 0.426278933;
cosLookup[11791] <= 0.426192199;
cosLookup[11792] <= 0.426105461;
cosLookup[11793] <= 0.426018719;
cosLookup[11794] <= 0.425931973;
cosLookup[11795] <= 0.425845224;
cosLookup[11796] <= 0.42575847;
cosLookup[11797] <= 0.425671713;
cosLookup[11798] <= 0.425584952;
cosLookup[11799] <= 0.425498186;
cosLookup[11800] <= 0.425411417;
cosLookup[11801] <= 0.425324644;
cosLookup[11802] <= 0.425237867;
cosLookup[11803] <= 0.425151086;
cosLookup[11804] <= 0.425064302;
cosLookup[11805] <= 0.424977513;
cosLookup[11806] <= 0.42489072;
cosLookup[11807] <= 0.424803924;
cosLookup[11808] <= 0.424717123;
cosLookup[11809] <= 0.424630319;
cosLookup[11810] <= 0.424543511;
cosLookup[11811] <= 0.424456699;
cosLookup[11812] <= 0.424369883;
cosLookup[11813] <= 0.424283063;
cosLookup[11814] <= 0.424196239;
cosLookup[11815] <= 0.424109411;
cosLookup[11816] <= 0.42402258;
cosLookup[11817] <= 0.423935744;
cosLookup[11818] <= 0.423848905;
cosLookup[11819] <= 0.423762062;
cosLookup[11820] <= 0.423675214;
cosLookup[11821] <= 0.423588363;
cosLookup[11822] <= 0.423501508;
cosLookup[11823] <= 0.423414649;
cosLookup[11824] <= 0.423327787;
cosLookup[11825] <= 0.42324092;
cosLookup[11826] <= 0.423154049;
cosLookup[11827] <= 0.423067175;
cosLookup[11828] <= 0.422980297;
cosLookup[11829] <= 0.422893414;
cosLookup[11830] <= 0.422806528;
cosLookup[11831] <= 0.422719638;
cosLookup[11832] <= 0.422632744;
cosLookup[11833] <= 0.422545847;
cosLookup[11834] <= 0.422458945;
cosLookup[11835] <= 0.422372039;
cosLookup[11836] <= 0.42228513;
cosLookup[11837] <= 0.422198217;
cosLookup[11838] <= 0.4221113;
cosLookup[11839] <= 0.422024379;
cosLookup[11840] <= 0.421937454;
cosLookup[11841] <= 0.421850525;
cosLookup[11842] <= 0.421763592;
cosLookup[11843] <= 0.421676655;
cosLookup[11844] <= 0.421589715;
cosLookup[11845] <= 0.421502771;
cosLookup[11846] <= 0.421415822;
cosLookup[11847] <= 0.42132887;
cosLookup[11848] <= 0.421241914;
cosLookup[11849] <= 0.421154955;
cosLookup[11850] <= 0.421067991;
cosLookup[11851] <= 0.420981023;
cosLookup[11852] <= 0.420894052;
cosLookup[11853] <= 0.420807077;
cosLookup[11854] <= 0.420720097;
cosLookup[11855] <= 0.420633114;
cosLookup[11856] <= 0.420546127;
cosLookup[11857] <= 0.420459137;
cosLookup[11858] <= 0.420372142;
cosLookup[11859] <= 0.420285144;
cosLookup[11860] <= 0.420198141;
cosLookup[11861] <= 0.420111135;
cosLookup[11862] <= 0.420024125;
cosLookup[11863] <= 0.419937111;
cosLookup[11864] <= 0.419850093;
cosLookup[11865] <= 0.419763071;
cosLookup[11866] <= 0.419676046;
cosLookup[11867] <= 0.419589016;
cosLookup[11868] <= 0.419501983;
cosLookup[11869] <= 0.419414946;
cosLookup[11870] <= 0.419327905;
cosLookup[11871] <= 0.41924086;
cosLookup[11872] <= 0.419153812;
cosLookup[11873] <= 0.419066759;
cosLookup[11874] <= 0.418979703;
cosLookup[11875] <= 0.418892643;
cosLookup[11876] <= 0.418805578;
cosLookup[11877] <= 0.418718511;
cosLookup[11878] <= 0.418631439;
cosLookup[11879] <= 0.418544363;
cosLookup[11880] <= 0.418457284;
cosLookup[11881] <= 0.4183702;
cosLookup[11882] <= 0.418283113;
cosLookup[11883] <= 0.418196022;
cosLookup[11884] <= 0.418108927;
cosLookup[11885] <= 0.418021829;
cosLookup[11886] <= 0.417934726;
cosLookup[11887] <= 0.41784762;
cosLookup[11888] <= 0.417760509;
cosLookup[11889] <= 0.417673395;
cosLookup[11890] <= 0.417586278;
cosLookup[11891] <= 0.417499156;
cosLookup[11892] <= 0.41741203;
cosLookup[11893] <= 0.417324901;
cosLookup[11894] <= 0.417237768;
cosLookup[11895] <= 0.41715063;
cosLookup[11896] <= 0.417063489;
cosLookup[11897] <= 0.416976345;
cosLookup[11898] <= 0.416889196;
cosLookup[11899] <= 0.416802044;
cosLookup[11900] <= 0.416714887;
cosLookup[11901] <= 0.416627727;
cosLookup[11902] <= 0.416540563;
cosLookup[11903] <= 0.416453396;
cosLookup[11904] <= 0.416366224;
cosLookup[11905] <= 0.416279049;
cosLookup[11906] <= 0.416191869;
cosLookup[11907] <= 0.416104686;
cosLookup[11908] <= 0.4160175;
cosLookup[11909] <= 0.415930309;
cosLookup[11910] <= 0.415843114;
cosLookup[11911] <= 0.415755916;
cosLookup[11912] <= 0.415668714;
cosLookup[11913] <= 0.415581508;
cosLookup[11914] <= 0.415494298;
cosLookup[11915] <= 0.415407084;
cosLookup[11916] <= 0.415319867;
cosLookup[11917] <= 0.415232646;
cosLookup[11918] <= 0.415145421;
cosLookup[11919] <= 0.415058192;
cosLookup[11920] <= 0.414970959;
cosLookup[11921] <= 0.414883722;
cosLookup[11922] <= 0.414796482;
cosLookup[11923] <= 0.414709238;
cosLookup[11924] <= 0.41462199;
cosLookup[11925] <= 0.414534738;
cosLookup[11926] <= 0.414447482;
cosLookup[11927] <= 0.414360223;
cosLookup[11928] <= 0.41427296;
cosLookup[11929] <= 0.414185693;
cosLookup[11930] <= 0.414098422;
cosLookup[11931] <= 0.414011147;
cosLookup[11932] <= 0.413923869;
cosLookup[11933] <= 0.413836587;
cosLookup[11934] <= 0.413749301;
cosLookup[11935] <= 0.413662011;
cosLookup[11936] <= 0.413574717;
cosLookup[11937] <= 0.41348742;
cosLookup[11938] <= 0.413400118;
cosLookup[11939] <= 0.413312813;
cosLookup[11940] <= 0.413225504;
cosLookup[11941] <= 0.413138192;
cosLookup[11942] <= 0.413050875;
cosLookup[11943] <= 0.412963555;
cosLookup[11944] <= 0.412876231;
cosLookup[11945] <= 0.412788903;
cosLookup[11946] <= 0.412701571;
cosLookup[11947] <= 0.412614236;
cosLookup[11948] <= 0.412526897;
cosLookup[11949] <= 0.412439554;
cosLookup[11950] <= 0.412352207;
cosLookup[11951] <= 0.412264856;
cosLookup[11952] <= 0.412177502;
cosLookup[11953] <= 0.412090144;
cosLookup[11954] <= 0.412002782;
cosLookup[11955] <= 0.411915416;
cosLookup[11956] <= 0.411828046;
cosLookup[11957] <= 0.411740673;
cosLookup[11958] <= 0.411653296;
cosLookup[11959] <= 0.411565915;
cosLookup[11960] <= 0.41147853;
cosLookup[11961] <= 0.411391142;
cosLookup[11962] <= 0.41130375;
cosLookup[11963] <= 0.411216354;
cosLookup[11964] <= 0.411128954;
cosLookup[11965] <= 0.41104155;
cosLookup[11966] <= 0.410954143;
cosLookup[11967] <= 0.410866732;
cosLookup[11968] <= 0.410779317;
cosLookup[11969] <= 0.410691898;
cosLookup[11970] <= 0.410604476;
cosLookup[11971] <= 0.410517049;
cosLookup[11972] <= 0.410429619;
cosLookup[11973] <= 0.410342186;
cosLookup[11974] <= 0.410254748;
cosLookup[11975] <= 0.410167307;
cosLookup[11976] <= 0.410079862;
cosLookup[11977] <= 0.409992413;
cosLookup[11978] <= 0.40990496;
cosLookup[11979] <= 0.409817504;
cosLookup[11980] <= 0.409730043;
cosLookup[11981] <= 0.409642579;
cosLookup[11982] <= 0.409555112;
cosLookup[11983] <= 0.40946764;
cosLookup[11984] <= 0.409380165;
cosLookup[11985] <= 0.409292686;
cosLookup[11986] <= 0.409205203;
cosLookup[11987] <= 0.409117717;
cosLookup[11988] <= 0.409030226;
cosLookup[11989] <= 0.408942732;
cosLookup[11990] <= 0.408855234;
cosLookup[11991] <= 0.408767733;
cosLookup[11992] <= 0.408680228;
cosLookup[11993] <= 0.408592718;
cosLookup[11994] <= 0.408505206;
cosLookup[11995] <= 0.408417689;
cosLookup[11996] <= 0.408330169;
cosLookup[11997] <= 0.408242645;
cosLookup[11998] <= 0.408155117;
cosLookup[11999] <= 0.408067585;
cosLookup[12000] <= 0.40798005;
cosLookup[12001] <= 0.407892511;
cosLookup[12002] <= 0.407804968;
cosLookup[12003] <= 0.407717421;
cosLookup[12004] <= 0.407629871;
cosLookup[12005] <= 0.407542317;
cosLookup[12006] <= 0.407454759;
cosLookup[12007] <= 0.407367197;
cosLookup[12008] <= 0.407279632;
cosLookup[12009] <= 0.407192063;
cosLookup[12010] <= 0.40710449;
cosLookup[12011] <= 0.407016913;
cosLookup[12012] <= 0.406929333;
cosLookup[12013] <= 0.406841749;
cosLookup[12014] <= 0.406754161;
cosLookup[12015] <= 0.40666657;
cosLookup[12016] <= 0.406578974;
cosLookup[12017] <= 0.406491375;
cosLookup[12018] <= 0.406403772;
cosLookup[12019] <= 0.406316166;
cosLookup[12020] <= 0.406228556;
cosLookup[12021] <= 0.406140942;
cosLookup[12022] <= 0.406053324;
cosLookup[12023] <= 0.405965703;
cosLookup[12024] <= 0.405878078;
cosLookup[12025] <= 0.405790449;
cosLookup[12026] <= 0.405702816;
cosLookup[12027] <= 0.40561518;
cosLookup[12028] <= 0.40552754;
cosLookup[12029] <= 0.405439896;
cosLookup[12030] <= 0.405352248;
cosLookup[12031] <= 0.405264597;
cosLookup[12032] <= 0.405176942;
cosLookup[12033] <= 0.405089283;
cosLookup[12034] <= 0.405001621;
cosLookup[12035] <= 0.404913955;
cosLookup[12036] <= 0.404826285;
cosLookup[12037] <= 0.404738611;
cosLookup[12038] <= 0.404650934;
cosLookup[12039] <= 0.404563253;
cosLookup[12040] <= 0.404475568;
cosLookup[12041] <= 0.40438788;
cosLookup[12042] <= 0.404300187;
cosLookup[12043] <= 0.404212492;
cosLookup[12044] <= 0.404124792;
cosLookup[12045] <= 0.404037089;
cosLookup[12046] <= 0.403949381;
cosLookup[12047] <= 0.403861671;
cosLookup[12048] <= 0.403773956;
cosLookup[12049] <= 0.403686238;
cosLookup[12050] <= 0.403598516;
cosLookup[12051] <= 0.40351079;
cosLookup[12052] <= 0.403423061;
cosLookup[12053] <= 0.403335328;
cosLookup[12054] <= 0.403247591;
cosLookup[12055] <= 0.403159851;
cosLookup[12056] <= 0.403072107;
cosLookup[12057] <= 0.402984359;
cosLookup[12058] <= 0.402896607;
cosLookup[12059] <= 0.402808852;
cosLookup[12060] <= 0.402721093;
cosLookup[12061] <= 0.40263333;
cosLookup[12062] <= 0.402545564;
cosLookup[12063] <= 0.402457794;
cosLookup[12064] <= 0.40237002;
cosLookup[12065] <= 0.402282243;
cosLookup[12066] <= 0.402194462;
cosLookup[12067] <= 0.402106677;
cosLookup[12068] <= 0.402018888;
cosLookup[12069] <= 0.401931096;
cosLookup[12070] <= 0.4018433;
cosLookup[12071] <= 0.4017555;
cosLookup[12072] <= 0.401667697;
cosLookup[12073] <= 0.40157989;
cosLookup[12074] <= 0.401492079;
cosLookup[12075] <= 0.401404265;
cosLookup[12076] <= 0.401316447;
cosLookup[12077] <= 0.401228625;
cosLookup[12078] <= 0.401140799;
cosLookup[12079] <= 0.40105297;
cosLookup[12080] <= 0.400965137;
cosLookup[12081] <= 0.400877301;
cosLookup[12082] <= 0.40078946;
cosLookup[12083] <= 0.400701617;
cosLookup[12084] <= 0.400613769;
cosLookup[12085] <= 0.400525918;
cosLookup[12086] <= 0.400438063;
cosLookup[12087] <= 0.400350204;
cosLookup[12088] <= 0.400262342;
cosLookup[12089] <= 0.400174476;
cosLookup[12090] <= 0.400086606;
cosLookup[12091] <= 0.399998733;
cosLookup[12092] <= 0.399910856;
cosLookup[12093] <= 0.399822975;
cosLookup[12094] <= 0.39973509;
cosLookup[12095] <= 0.399647202;
cosLookup[12096] <= 0.399559311;
cosLookup[12097] <= 0.399471415;
cosLookup[12098] <= 0.399383516;
cosLookup[12099] <= 0.399295613;
cosLookup[12100] <= 0.399207707;
cosLookup[12101] <= 0.399119797;
cosLookup[12102] <= 0.399031883;
cosLookup[12103] <= 0.398943966;
cosLookup[12104] <= 0.398856045;
cosLookup[12105] <= 0.39876812;
cosLookup[12106] <= 0.398680191;
cosLookup[12107] <= 0.398592259;
cosLookup[12108] <= 0.398504323;
cosLookup[12109] <= 0.398416384;
cosLookup[12110] <= 0.398328441;
cosLookup[12111] <= 0.398240494;
cosLookup[12112] <= 0.398152544;
cosLookup[12113] <= 0.39806459;
cosLookup[12114] <= 0.397976632;
cosLookup[12115] <= 0.397888671;
cosLookup[12116] <= 0.397800706;
cosLookup[12117] <= 0.397712737;
cosLookup[12118] <= 0.397624764;
cosLookup[12119] <= 0.397536788;
cosLookup[12120] <= 0.397448809;
cosLookup[12121] <= 0.397360825;
cosLookup[12122] <= 0.397272838;
cosLookup[12123] <= 0.397184848;
cosLookup[12124] <= 0.397096854;
cosLookup[12125] <= 0.397008856;
cosLookup[12126] <= 0.396920854;
cosLookup[12127] <= 0.396832849;
cosLookup[12128] <= 0.39674484;
cosLookup[12129] <= 0.396656827;
cosLookup[12130] <= 0.396568811;
cosLookup[12131] <= 0.396480791;
cosLookup[12132] <= 0.396392768;
cosLookup[12133] <= 0.396304741;
cosLookup[12134] <= 0.39621671;
cosLookup[12135] <= 0.396128676;
cosLookup[12136] <= 0.396040638;
cosLookup[12137] <= 0.395952596;
cosLookup[12138] <= 0.395864551;
cosLookup[12139] <= 0.395776502;
cosLookup[12140] <= 0.395688449;
cosLookup[12141] <= 0.395600393;
cosLookup[12142] <= 0.395512333;
cosLookup[12143] <= 0.395424269;
cosLookup[12144] <= 0.395336202;
cosLookup[12145] <= 0.395248131;
cosLookup[12146] <= 0.395160057;
cosLookup[12147] <= 0.395071979;
cosLookup[12148] <= 0.394983897;
cosLookup[12149] <= 0.394895812;
cosLookup[12150] <= 0.394807723;
cosLookup[12151] <= 0.394719631;
cosLookup[12152] <= 0.394631534;
cosLookup[12153] <= 0.394543435;
cosLookup[12154] <= 0.394455331;
cosLookup[12155] <= 0.394367224;
cosLookup[12156] <= 0.394279113;
cosLookup[12157] <= 0.394190999;
cosLookup[12158] <= 0.394102881;
cosLookup[12159] <= 0.394014759;
cosLookup[12160] <= 0.393926634;
cosLookup[12161] <= 0.393838505;
cosLookup[12162] <= 0.393750373;
cosLookup[12163] <= 0.393662237;
cosLookup[12164] <= 0.393574097;
cosLookup[12165] <= 0.393485954;
cosLookup[12166] <= 0.393397807;
cosLookup[12167] <= 0.393309657;
cosLookup[12168] <= 0.393221502;
cosLookup[12169] <= 0.393133345;
cosLookup[12170] <= 0.393045183;
cosLookup[12171] <= 0.392957018;
cosLookup[12172] <= 0.39286885;
cosLookup[12173] <= 0.392780678;
cosLookup[12174] <= 0.392692502;
cosLookup[12175] <= 0.392604322;
cosLookup[12176] <= 0.392516139;
cosLookup[12177] <= 0.392427953;
cosLookup[12178] <= 0.392339762;
cosLookup[12179] <= 0.392251569;
cosLookup[12180] <= 0.392163371;
cosLookup[12181] <= 0.39207517;
cosLookup[12182] <= 0.391986965;
cosLookup[12183] <= 0.391898757;
cosLookup[12184] <= 0.391810545;
cosLookup[12185] <= 0.39172233;
cosLookup[12186] <= 0.391634111;
cosLookup[12187] <= 0.391545888;
cosLookup[12188] <= 0.391457662;
cosLookup[12189] <= 0.391369432;
cosLookup[12190] <= 0.391281198;
cosLookup[12191] <= 0.391192961;
cosLookup[12192] <= 0.39110472;
cosLookup[12193] <= 0.391016476;
cosLookup[12194] <= 0.390928228;
cosLookup[12195] <= 0.390839977;
cosLookup[12196] <= 0.390751722;
cosLookup[12197] <= 0.390663463;
cosLookup[12198] <= 0.390575201;
cosLookup[12199] <= 0.390486935;
cosLookup[12200] <= 0.390398666;
cosLookup[12201] <= 0.390310393;
cosLookup[12202] <= 0.390222116;
cosLookup[12203] <= 0.390133836;
cosLookup[12204] <= 0.390045552;
cosLookup[12205] <= 0.389957265;
cosLookup[12206] <= 0.389868974;
cosLookup[12207] <= 0.389780679;
cosLookup[12208] <= 0.389692381;
cosLookup[12209] <= 0.38960408;
cosLookup[12210] <= 0.389515774;
cosLookup[12211] <= 0.389427465;
cosLookup[12212] <= 0.389339153;
cosLookup[12213] <= 0.389250837;
cosLookup[12214] <= 0.389162517;
cosLookup[12215] <= 0.389074194;
cosLookup[12216] <= 0.388985868;
cosLookup[12217] <= 0.388897537;
cosLookup[12218] <= 0.388809203;
cosLookup[12219] <= 0.388720866;
cosLookup[12220] <= 0.388632525;
cosLookup[12221] <= 0.38854418;
cosLookup[12222] <= 0.388455832;
cosLookup[12223] <= 0.38836748;
cosLookup[12224] <= 0.388279125;
cosLookup[12225] <= 0.388190766;
cosLookup[12226] <= 0.388102404;
cosLookup[12227] <= 0.388014038;
cosLookup[12228] <= 0.387925668;
cosLookup[12229] <= 0.387837295;
cosLookup[12230] <= 0.387748918;
cosLookup[12231] <= 0.387660538;
cosLookup[12232] <= 0.387572154;
cosLookup[12233] <= 0.387483767;
cosLookup[12234] <= 0.387395376;
cosLookup[12235] <= 0.387306981;
cosLookup[12236] <= 0.387218583;
cosLookup[12237] <= 0.387130181;
cosLookup[12238] <= 0.387041776;
cosLookup[12239] <= 0.386953367;
cosLookup[12240] <= 0.386864955;
cosLookup[12241] <= 0.386776539;
cosLookup[12242] <= 0.38668812;
cosLookup[12243] <= 0.386599697;
cosLookup[12244] <= 0.38651127;
cosLookup[12245] <= 0.38642284;
cosLookup[12246] <= 0.386334406;
cosLookup[12247] <= 0.386245969;
cosLookup[12248] <= 0.386157528;
cosLookup[12249] <= 0.386069084;
cosLookup[12250] <= 0.385980636;
cosLookup[12251] <= 0.385892185;
cosLookup[12252] <= 0.38580373;
cosLookup[12253] <= 0.385715271;
cosLookup[12254] <= 0.385626809;
cosLookup[12255] <= 0.385538344;
cosLookup[12256] <= 0.385449874;
cosLookup[12257] <= 0.385361402;
cosLookup[12258] <= 0.385272926;
cosLookup[12259] <= 0.385184446;
cosLookup[12260] <= 0.385095962;
cosLookup[12261] <= 0.385007476;
cosLookup[12262] <= 0.384918985;
cosLookup[12263] <= 0.384830491;
cosLookup[12264] <= 0.384741994;
cosLookup[12265] <= 0.384653493;
cosLookup[12266] <= 0.384564988;
cosLookup[12267] <= 0.38447648;
cosLookup[12268] <= 0.384387969;
cosLookup[12269] <= 0.384299453;
cosLookup[12270] <= 0.384210935;
cosLookup[12271] <= 0.384122413;
cosLookup[12272] <= 0.384033887;
cosLookup[12273] <= 0.383945358;
cosLookup[12274] <= 0.383856825;
cosLookup[12275] <= 0.383768288;
cosLookup[12276] <= 0.383679749;
cosLookup[12277] <= 0.383591205;
cosLookup[12278] <= 0.383502658;
cosLookup[12279] <= 0.383414108;
cosLookup[12280] <= 0.383325554;
cosLookup[12281] <= 0.383236996;
cosLookup[12282] <= 0.383148435;
cosLookup[12283] <= 0.383059871;
cosLookup[12284] <= 0.382971303;
cosLookup[12285] <= 0.382882731;
cosLookup[12286] <= 0.382794156;
cosLookup[12287] <= 0.382705578;
cosLookup[12288] <= 0.382616995;
cosLookup[12289] <= 0.38252841;
cosLookup[12290] <= 0.382439821;
cosLookup[12291] <= 0.382351228;
cosLookup[12292] <= 0.382262632;
cosLookup[12293] <= 0.382174032;
cosLookup[12294] <= 0.382085429;
cosLookup[12295] <= 0.381996822;
cosLookup[12296] <= 0.381908212;
cosLookup[12297] <= 0.381819598;
cosLookup[12298] <= 0.381730981;
cosLookup[12299] <= 0.38164236;
cosLookup[12300] <= 0.381553736;
cosLookup[12301] <= 0.381465108;
cosLookup[12302] <= 0.381376477;
cosLookup[12303] <= 0.381287842;
cosLookup[12304] <= 0.381199204;
cosLookup[12305] <= 0.381110562;
cosLookup[12306] <= 0.381021916;
cosLookup[12307] <= 0.380933268;
cosLookup[12308] <= 0.380844615;
cosLookup[12309] <= 0.38075596;
cosLookup[12310] <= 0.3806673;
cosLookup[12311] <= 0.380578637;
cosLookup[12312] <= 0.380489971;
cosLookup[12313] <= 0.380401301;
cosLookup[12314] <= 0.380312628;
cosLookup[12315] <= 0.380223951;
cosLookup[12316] <= 0.380135271;
cosLookup[12317] <= 0.380046587;
cosLookup[12318] <= 0.3799579;
cosLookup[12319] <= 0.379869209;
cosLookup[12320] <= 0.379780515;
cosLookup[12321] <= 0.379691817;
cosLookup[12322] <= 0.379603116;
cosLookup[12323] <= 0.379514411;
cosLookup[12324] <= 0.379425703;
cosLookup[12325] <= 0.379336991;
cosLookup[12326] <= 0.379248276;
cosLookup[12327] <= 0.379159557;
cosLookup[12328] <= 0.379070835;
cosLookup[12329] <= 0.378982109;
cosLookup[12330] <= 0.37889338;
cosLookup[12331] <= 0.378804647;
cosLookup[12332] <= 0.378715911;
cosLookup[12333] <= 0.378627172;
cosLookup[12334] <= 0.378538429;
cosLookup[12335] <= 0.378449682;
cosLookup[12336] <= 0.378360932;
cosLookup[12337] <= 0.378272178;
cosLookup[12338] <= 0.378183421;
cosLookup[12339] <= 0.378094661;
cosLookup[12340] <= 0.378005897;
cosLookup[12341] <= 0.37791713;
cosLookup[12342] <= 0.377828359;
cosLookup[12343] <= 0.377739584;
cosLookup[12344] <= 0.377650806;
cosLookup[12345] <= 0.377562025;
cosLookup[12346] <= 0.37747324;
cosLookup[12347] <= 0.377384452;
cosLookup[12348] <= 0.37729566;
cosLookup[12349] <= 0.377206865;
cosLookup[12350] <= 0.377118067;
cosLookup[12351] <= 0.377029264;
cosLookup[12352] <= 0.376940459;
cosLookup[12353] <= 0.37685165;
cosLookup[12354] <= 0.376762837;
cosLookup[12355] <= 0.376674021;
cosLookup[12356] <= 0.376585202;
cosLookup[12357] <= 0.376496379;
cosLookup[12358] <= 0.376407552;
cosLookup[12359] <= 0.376318723;
cosLookup[12360] <= 0.376229889;
cosLookup[12361] <= 0.376141053;
cosLookup[12362] <= 0.376052212;
cosLookup[12363] <= 0.375963369;
cosLookup[12364] <= 0.375874522;
cosLookup[12365] <= 0.375785671;
cosLookup[12366] <= 0.375696817;
cosLookup[12367] <= 0.37560796;
cosLookup[12368] <= 0.375519099;
cosLookup[12369] <= 0.375430234;
cosLookup[12370] <= 0.375341366;
cosLookup[12371] <= 0.375252495;
cosLookup[12372] <= 0.37516362;
cosLookup[12373] <= 0.375074742;
cosLookup[12374] <= 0.37498586;
cosLookup[12375] <= 0.374896975;
cosLookup[12376] <= 0.374808087;
cosLookup[12377] <= 0.374719195;
cosLookup[12378] <= 0.374630299;
cosLookup[12379] <= 0.374541401;
cosLookup[12380] <= 0.374452498;
cosLookup[12381] <= 0.374363593;
cosLookup[12382] <= 0.374274683;
cosLookup[12383] <= 0.374185771;
cosLookup[12384] <= 0.374096855;
cosLookup[12385] <= 0.374007935;
cosLookup[12386] <= 0.373919012;
cosLookup[12387] <= 0.373830086;
cosLookup[12388] <= 0.373741156;
cosLookup[12389] <= 0.373652223;
cosLookup[12390] <= 0.373563286;
cosLookup[12391] <= 0.373474346;
cosLookup[12392] <= 0.373385402;
cosLookup[12393] <= 0.373296455;
cosLookup[12394] <= 0.373207505;
cosLookup[12395] <= 0.373118551;
cosLookup[12396] <= 0.373029594;
cosLookup[12397] <= 0.372940633;
cosLookup[12398] <= 0.372851669;
cosLookup[12399] <= 0.372762701;
cosLookup[12400] <= 0.37267373;
cosLookup[12401] <= 0.372584756;
cosLookup[12402] <= 0.372495778;
cosLookup[12403] <= 0.372406797;
cosLookup[12404] <= 0.372317812;
cosLookup[12405] <= 0.372228824;
cosLookup[12406] <= 0.372139832;
cosLookup[12407] <= 0.372050837;
cosLookup[12408] <= 0.371961839;
cosLookup[12409] <= 0.371872837;
cosLookup[12410] <= 0.371783832;
cosLookup[12411] <= 0.371694823;
cosLookup[12412] <= 0.371605811;
cosLookup[12413] <= 0.371516796;
cosLookup[12414] <= 0.371427777;
cosLookup[12415] <= 0.371338755;
cosLookup[12416] <= 0.371249729;
cosLookup[12417] <= 0.3711607;
cosLookup[12418] <= 0.371071667;
cosLookup[12419] <= 0.370982631;
cosLookup[12420] <= 0.370893592;
cosLookup[12421] <= 0.370804549;
cosLookup[12422] <= 0.370715503;
cosLookup[12423] <= 0.370626453;
cosLookup[12424] <= 0.3705374;
cosLookup[12425] <= 0.370448344;
cosLookup[12426] <= 0.370359284;
cosLookup[12427] <= 0.370270221;
cosLookup[12428] <= 0.370181154;
cosLookup[12429] <= 0.370092084;
cosLookup[12430] <= 0.370003011;
cosLookup[12431] <= 0.369913934;
cosLookup[12432] <= 0.369824854;
cosLookup[12433] <= 0.36973577;
cosLookup[12434] <= 0.369646683;
cosLookup[12435] <= 0.369557593;
cosLookup[12436] <= 0.369468499;
cosLookup[12437] <= 0.369379402;
cosLookup[12438] <= 0.369290301;
cosLookup[12439] <= 0.369201197;
cosLookup[12440] <= 0.36911209;
cosLookup[12441] <= 0.369022979;
cosLookup[12442] <= 0.368933865;
cosLookup[12443] <= 0.368844747;
cosLookup[12444] <= 0.368755626;
cosLookup[12445] <= 0.368666502;
cosLookup[12446] <= 0.368577374;
cosLookup[12447] <= 0.368488243;
cosLookup[12448] <= 0.368399108;
cosLookup[12449] <= 0.36830997;
cosLookup[12450] <= 0.368220829;
cosLookup[12451] <= 0.368131684;
cosLookup[12452] <= 0.368042536;
cosLookup[12453] <= 0.367953385;
cosLookup[12454] <= 0.36786423;
cosLookup[12455] <= 0.367775072;
cosLookup[12456] <= 0.36768591;
cosLookup[12457] <= 0.367596745;
cosLookup[12458] <= 0.367507577;
cosLookup[12459] <= 0.367418405;
cosLookup[12460] <= 0.36732923;
cosLookup[12461] <= 0.367240052;
cosLookup[12462] <= 0.36715087;
cosLookup[12463] <= 0.367061684;
cosLookup[12464] <= 0.366972496;
cosLookup[12465] <= 0.366883304;
cosLookup[12466] <= 0.366794109;
cosLookup[12467] <= 0.36670491;
cosLookup[12468] <= 0.366615708;
cosLookup[12469] <= 0.366526502;
cosLookup[12470] <= 0.366437293;
cosLookup[12471] <= 0.366348081;
cosLookup[12472] <= 0.366258866;
cosLookup[12473] <= 0.366169647;
cosLookup[12474] <= 0.366080424;
cosLookup[12475] <= 0.365991199;
cosLookup[12476] <= 0.36590197;
cosLookup[12477] <= 0.365812737;
cosLookup[12478] <= 0.365723501;
cosLookup[12479] <= 0.365634262;
cosLookup[12480] <= 0.36554502;
cosLookup[12481] <= 0.365455774;
cosLookup[12482] <= 0.365366525;
cosLookup[12483] <= 0.365277272;
cosLookup[12484] <= 0.365188016;
cosLookup[12485] <= 0.365098757;
cosLookup[12486] <= 0.365009494;
cosLookup[12487] <= 0.364920228;
cosLookup[12488] <= 0.364830959;
cosLookup[12489] <= 0.364741686;
cosLookup[12490] <= 0.36465241;
cosLookup[12491] <= 0.364563131;
cosLookup[12492] <= 0.364473848;
cosLookup[12493] <= 0.364384562;
cosLookup[12494] <= 0.364295272;
cosLookup[12495] <= 0.36420598;
cosLookup[12496] <= 0.364116684;
cosLookup[12497] <= 0.364027384;
cosLookup[12498] <= 0.363938081;
cosLookup[12499] <= 0.363848775;
cosLookup[12500] <= 0.363759465;
cosLookup[12501] <= 0.363670153;
cosLookup[12502] <= 0.363580836;
cosLookup[12503] <= 0.363491517;
cosLookup[12504] <= 0.363402194;
cosLookup[12505] <= 0.363312868;
cosLookup[12506] <= 0.363223538;
cosLookup[12507] <= 0.363134205;
cosLookup[12508] <= 0.363044869;
cosLookup[12509] <= 0.362955529;
cosLookup[12510] <= 0.362866186;
cosLookup[12511] <= 0.36277684;
cosLookup[12512] <= 0.36268749;
cosLookup[12513] <= 0.362598137;
cosLookup[12514] <= 0.362508781;
cosLookup[12515] <= 0.362419421;
cosLookup[12516] <= 0.362330058;
cosLookup[12517] <= 0.362240692;
cosLookup[12518] <= 0.362151323;
cosLookup[12519] <= 0.36206195;
cosLookup[12520] <= 0.361972573;
cosLookup[12521] <= 0.361883194;
cosLookup[12522] <= 0.361793811;
cosLookup[12523] <= 0.361704425;
cosLookup[12524] <= 0.361615035;
cosLookup[12525] <= 0.361525642;
cosLookup[12526] <= 0.361436246;
cosLookup[12527] <= 0.361346846;
cosLookup[12528] <= 0.361257444;
cosLookup[12529] <= 0.361168037;
cosLookup[12530] <= 0.361078628;
cosLookup[12531] <= 0.360989215;
cosLookup[12532] <= 0.360899799;
cosLookup[12533] <= 0.360810379;
cosLookup[12534] <= 0.360720957;
cosLookup[12535] <= 0.360631531;
cosLookup[12536] <= 0.360542101;
cosLookup[12537] <= 0.360452668;
cosLookup[12538] <= 0.360363232;
cosLookup[12539] <= 0.360273793;
cosLookup[12540] <= 0.36018435;
cosLookup[12541] <= 0.360094904;
cosLookup[12542] <= 0.360005455;
cosLookup[12543] <= 0.359916002;
cosLookup[12544] <= 0.359826547;
cosLookup[12545] <= 0.359737087;
cosLookup[12546] <= 0.359647625;
cosLookup[12547] <= 0.359558159;
cosLookup[12548] <= 0.35946869;
cosLookup[12549] <= 0.359379217;
cosLookup[12550] <= 0.359289742;
cosLookup[12551] <= 0.359200263;
cosLookup[12552] <= 0.35911078;
cosLookup[12553] <= 0.359021295;
cosLookup[12554] <= 0.358931806;
cosLookup[12555] <= 0.358842313;
cosLookup[12556] <= 0.358752818;
cosLookup[12557] <= 0.358663319;
cosLookup[12558] <= 0.358573817;
cosLookup[12559] <= 0.358484312;
cosLookup[12560] <= 0.358394803;
cosLookup[12561] <= 0.358305291;
cosLookup[12562] <= 0.358215775;
cosLookup[12563] <= 0.358126257;
cosLookup[12564] <= 0.358036735;
cosLookup[12565] <= 0.35794721;
cosLookup[12566] <= 0.357857681;
cosLookup[12567] <= 0.357768149;
cosLookup[12568] <= 0.357678614;
cosLookup[12569] <= 0.357589076;
cosLookup[12570] <= 0.357499534;
cosLookup[12571] <= 0.35740999;
cosLookup[12572] <= 0.357320441;
cosLookup[12573] <= 0.35723089;
cosLookup[12574] <= 0.357141335;
cosLookup[12575] <= 0.357051777;
cosLookup[12576] <= 0.356962216;
cosLookup[12577] <= 0.356872651;
cosLookup[12578] <= 0.356783083;
cosLookup[12579] <= 0.356693512;
cosLookup[12580] <= 0.356603937;
cosLookup[12581] <= 0.35651436;
cosLookup[12582] <= 0.356424779;
cosLookup[12583] <= 0.356335194;
cosLookup[12584] <= 0.356245607;
cosLookup[12585] <= 0.356156016;
cosLookup[12586] <= 0.356066422;
cosLookup[12587] <= 0.355976824;
cosLookup[12588] <= 0.355887224;
cosLookup[12589] <= 0.35579762;
cosLookup[12590] <= 0.355708013;
cosLookup[12591] <= 0.355618402;
cosLookup[12592] <= 0.355528788;
cosLookup[12593] <= 0.355439171;
cosLookup[12594] <= 0.355349551;
cosLookup[12595] <= 0.355259927;
cosLookup[12596] <= 0.355170301;
cosLookup[12597] <= 0.355080671;
cosLookup[12598] <= 0.354991037;
cosLookup[12599] <= 0.354901401;
cosLookup[12600] <= 0.354811761;
cosLookup[12601] <= 0.354722118;
cosLookup[12602] <= 0.354632471;
cosLookup[12603] <= 0.354542822;
cosLookup[12604] <= 0.354453169;
cosLookup[12605] <= 0.354363512;
cosLookup[12606] <= 0.354273853;
cosLookup[12607] <= 0.35418419;
cosLookup[12608] <= 0.354094524;
cosLookup[12609] <= 0.354004855;
cosLookup[12610] <= 0.353915183;
cosLookup[12611] <= 0.353825507;
cosLookup[12612] <= 0.353735828;
cosLookup[12613] <= 0.353646146;
cosLookup[12614] <= 0.35355646;
cosLookup[12615] <= 0.353466772;
cosLookup[12616] <= 0.35337708;
cosLookup[12617] <= 0.353287384;
cosLookup[12618] <= 0.353197686;
cosLookup[12619] <= 0.353107984;
cosLookup[12620] <= 0.353018279;
cosLookup[12621] <= 0.352928571;
cosLookup[12622] <= 0.35283886;
cosLookup[12623] <= 0.352749145;
cosLookup[12624] <= 0.352659427;
cosLookup[12625] <= 0.352569706;
cosLookup[12626] <= 0.352479982;
cosLookup[12627] <= 0.352390254;
cosLookup[12628] <= 0.352300523;
cosLookup[12629] <= 0.352210789;
cosLookup[12630] <= 0.352121051;
cosLookup[12631] <= 0.352031311;
cosLookup[12632] <= 0.351941567;
cosLookup[12633] <= 0.35185182;
cosLookup[12634] <= 0.35176207;
cosLookup[12635] <= 0.351672316;
cosLookup[12636] <= 0.351582559;
cosLookup[12637] <= 0.351492799;
cosLookup[12638] <= 0.351403036;
cosLookup[12639] <= 0.35131327;
cosLookup[12640] <= 0.3512235;
cosLookup[12641] <= 0.351133727;
cosLookup[12642] <= 0.351043951;
cosLookup[12643] <= 0.350954171;
cosLookup[12644] <= 0.350864389;
cosLookup[12645] <= 0.350774603;
cosLookup[12646] <= 0.350684814;
cosLookup[12647] <= 0.350595022;
cosLookup[12648] <= 0.350505226;
cosLookup[12649] <= 0.350415427;
cosLookup[12650] <= 0.350325625;
cosLookup[12651] <= 0.35023582;
cosLookup[12652] <= 0.350146012;
cosLookup[12653] <= 0.3500562;
cosLookup[12654] <= 0.349966385;
cosLookup[12655] <= 0.349876567;
cosLookup[12656] <= 0.349786746;
cosLookup[12657] <= 0.349696922;
cosLookup[12658] <= 0.349607094;
cosLookup[12659] <= 0.349517263;
cosLookup[12660] <= 0.349427429;
cosLookup[12661] <= 0.349337592;
cosLookup[12662] <= 0.349247751;
cosLookup[12663] <= 0.349157907;
cosLookup[12664] <= 0.34906806;
cosLookup[12665] <= 0.34897821;
cosLookup[12666] <= 0.348888357;
cosLookup[12667] <= 0.3487985;
cosLookup[12668] <= 0.34870864;
cosLookup[12669] <= 0.348618777;
cosLookup[12670] <= 0.348528911;
cosLookup[12671] <= 0.348439042;
cosLookup[12672] <= 0.348349169;
cosLookup[12673] <= 0.348259293;
cosLookup[12674] <= 0.348169414;
cosLookup[12675] <= 0.348079532;
cosLookup[12676] <= 0.347989647;
cosLookup[12677] <= 0.347899758;
cosLookup[12678] <= 0.347809866;
cosLookup[12679] <= 0.347719971;
cosLookup[12680] <= 0.347630073;
cosLookup[12681] <= 0.347540172;
cosLookup[12682] <= 0.347450267;
cosLookup[12683] <= 0.347360359;
cosLookup[12684] <= 0.347270448;
cosLookup[12685] <= 0.347180534;
cosLookup[12686] <= 0.347090617;
cosLookup[12687] <= 0.347000696;
cosLookup[12688] <= 0.346910772;
cosLookup[12689] <= 0.346820845;
cosLookup[12690] <= 0.346730915;
cosLookup[12691] <= 0.346640982;
cosLookup[12692] <= 0.346551045;
cosLookup[12693] <= 0.346461106;
cosLookup[12694] <= 0.346371163;
cosLookup[12695] <= 0.346281217;
cosLookup[12696] <= 0.346191268;
cosLookup[12697] <= 0.346101315;
cosLookup[12698] <= 0.34601136;
cosLookup[12699] <= 0.345921401;
cosLookup[12700] <= 0.345831439;
cosLookup[12701] <= 0.345741474;
cosLookup[12702] <= 0.345651505;
cosLookup[12703] <= 0.345561534;
cosLookup[12704] <= 0.345471559;
cosLookup[12705] <= 0.345381581;
cosLookup[12706] <= 0.3452916;
cosLookup[12707] <= 0.345201616;
cosLookup[12708] <= 0.345111629;
cosLookup[12709] <= 0.345021638;
cosLookup[12710] <= 0.344931644;
cosLookup[12711] <= 0.344841648;
cosLookup[12712] <= 0.344751647;
cosLookup[12713] <= 0.344661644;
cosLookup[12714] <= 0.344571638;
cosLookup[12715] <= 0.344481628;
cosLookup[12716] <= 0.344391616;
cosLookup[12717] <= 0.3443016;
cosLookup[12718] <= 0.344211581;
cosLookup[12719] <= 0.344121558;
cosLookup[12720] <= 0.344031533;
cosLookup[12721] <= 0.343941504;
cosLookup[12722] <= 0.343851473;
cosLookup[12723] <= 0.343761438;
cosLookup[12724] <= 0.3436714;
cosLookup[12725] <= 0.343581359;
cosLookup[12726] <= 0.343491314;
cosLookup[12727] <= 0.343401267;
cosLookup[12728] <= 0.343311216;
cosLookup[12729] <= 0.343221162;
cosLookup[12730] <= 0.343131105;
cosLookup[12731] <= 0.343041045;
cosLookup[12732] <= 0.342950982;
cosLookup[12733] <= 0.342860915;
cosLookup[12734] <= 0.342770846;
cosLookup[12735] <= 0.342680773;
cosLookup[12736] <= 0.342590697;
cosLookup[12737] <= 0.342500618;
cosLookup[12738] <= 0.342410536;
cosLookup[12739] <= 0.342320451;
cosLookup[12740] <= 0.342230362;
cosLookup[12741] <= 0.34214027;
cosLookup[12742] <= 0.342050176;
cosLookup[12743] <= 0.341960078;
cosLookup[12744] <= 0.341869977;
cosLookup[12745] <= 0.341779872;
cosLookup[12746] <= 0.341689765;
cosLookup[12747] <= 0.341599655;
cosLookup[12748] <= 0.341509541;
cosLookup[12749] <= 0.341419424;
cosLookup[12750] <= 0.341329304;
cosLookup[12751] <= 0.341239181;
cosLookup[12752] <= 0.341149055;
cosLookup[12753] <= 0.341058926;
cosLookup[12754] <= 0.340968793;
cosLookup[12755] <= 0.340878658;
cosLookup[12756] <= 0.340788519;
cosLookup[12757] <= 0.340698377;
cosLookup[12758] <= 0.340608232;
cosLookup[12759] <= 0.340518084;
cosLookup[12760] <= 0.340427933;
cosLookup[12761] <= 0.340337778;
cosLookup[12762] <= 0.340247621;
cosLookup[12763] <= 0.34015746;
cosLookup[12764] <= 0.340067296;
cosLookup[12765] <= 0.339977129;
cosLookup[12766] <= 0.339886959;
cosLookup[12767] <= 0.339796786;
cosLookup[12768] <= 0.33970661;
cosLookup[12769] <= 0.339616431;
cosLookup[12770] <= 0.339526248;
cosLookup[12771] <= 0.339436063;
cosLookup[12772] <= 0.339345874;
cosLookup[12773] <= 0.339255682;
cosLookup[12774] <= 0.339165487;
cosLookup[12775] <= 0.339075289;
cosLookup[12776] <= 0.338985088;
cosLookup[12777] <= 0.338894883;
cosLookup[12778] <= 0.338804676;
cosLookup[12779] <= 0.338714465;
cosLookup[12780] <= 0.338624252;
cosLookup[12781] <= 0.338534035;
cosLookup[12782] <= 0.338443815;
cosLookup[12783] <= 0.338353592;
cosLookup[12784] <= 0.338263366;
cosLookup[12785] <= 0.338173136;
cosLookup[12786] <= 0.338082904;
cosLookup[12787] <= 0.337992669;
cosLookup[12788] <= 0.33790243;
cosLookup[12789] <= 0.337812188;
cosLookup[12790] <= 0.337721944;
cosLookup[12791] <= 0.337631696;
cosLookup[12792] <= 0.337541445;
cosLookup[12793] <= 0.337451191;
cosLookup[12794] <= 0.337360933;
cosLookup[12795] <= 0.337270673;
cosLookup[12796] <= 0.33718041;
cosLookup[12797] <= 0.337090143;
cosLookup[12798] <= 0.336999874;
cosLookup[12799] <= 0.336909601;
cosLookup[12800] <= 0.336819325;
cosLookup[12801] <= 0.336729046;
cosLookup[12802] <= 0.336638764;
cosLookup[12803] <= 0.336548479;
cosLookup[12804] <= 0.336458191;
cosLookup[12805] <= 0.3363679;
cosLookup[12806] <= 0.336277605;
cosLookup[12807] <= 0.336187308;
cosLookup[12808] <= 0.336097007;
cosLookup[12809] <= 0.336006704;
cosLookup[12810] <= 0.335916397;
cosLookup[12811] <= 0.335826087;
cosLookup[12812] <= 0.335735774;
cosLookup[12813] <= 0.335645458;
cosLookup[12814] <= 0.335555139;
cosLookup[12815] <= 0.335464817;
cosLookup[12816] <= 0.335374492;
cosLookup[12817] <= 0.335284164;
cosLookup[12818] <= 0.335193832;
cosLookup[12819] <= 0.335103498;
cosLookup[12820] <= 0.33501316;
cosLookup[12821] <= 0.33492282;
cosLookup[12822] <= 0.334832476;
cosLookup[12823] <= 0.334742129;
cosLookup[12824] <= 0.334651779;
cosLookup[12825] <= 0.334561426;
cosLookup[12826] <= 0.33447107;
cosLookup[12827] <= 0.334380711;
cosLookup[12828] <= 0.334290349;
cosLookup[12829] <= 0.334199984;
cosLookup[12830] <= 0.334109615;
cosLookup[12831] <= 0.334019244;
cosLookup[12832] <= 0.33392887;
cosLookup[12833] <= 0.333838492;
cosLookup[12834] <= 0.333748111;
cosLookup[12835] <= 0.333657728;
cosLookup[12836] <= 0.333567341;
cosLookup[12837] <= 0.333476951;
cosLookup[12838] <= 0.333386558;
cosLookup[12839] <= 0.333296163;
cosLookup[12840] <= 0.333205764;
cosLookup[12841] <= 0.333115361;
cosLookup[12842] <= 0.333024956;
cosLookup[12843] <= 0.332934548;
cosLookup[12844] <= 0.332844137;
cosLookup[12845] <= 0.332753723;
cosLookup[12846] <= 0.332663305;
cosLookup[12847] <= 0.332572885;
cosLookup[12848] <= 0.332482461;
cosLookup[12849] <= 0.332392035;
cosLookup[12850] <= 0.332301605;
cosLookup[12851] <= 0.332211173;
cosLookup[12852] <= 0.332120737;
cosLookup[12853] <= 0.332030298;
cosLookup[12854] <= 0.331939856;
cosLookup[12855] <= 0.331849411;
cosLookup[12856] <= 0.331758964;
cosLookup[12857] <= 0.331668513;
cosLookup[12858] <= 0.331578059;
cosLookup[12859] <= 0.331487602;
cosLookup[12860] <= 0.331397141;
cosLookup[12861] <= 0.331306678;
cosLookup[12862] <= 0.331216212;
cosLookup[12863] <= 0.331125743;
cosLookup[12864] <= 0.331035271;
cosLookup[12865] <= 0.330944795;
cosLookup[12866] <= 0.330854317;
cosLookup[12867] <= 0.330763836;
cosLookup[12868] <= 0.330673351;
cosLookup[12869] <= 0.330582864;
cosLookup[12870] <= 0.330492373;
cosLookup[12871] <= 0.33040188;
cosLookup[12872] <= 0.330311383;
cosLookup[12873] <= 0.330220883;
cosLookup[12874] <= 0.330130381;
cosLookup[12875] <= 0.330039875;
cosLookup[12876] <= 0.329949366;
cosLookup[12877] <= 0.329858854;
cosLookup[12878] <= 0.32976834;
cosLookup[12879] <= 0.329677822;
cosLookup[12880] <= 0.329587301;
cosLookup[12881] <= 0.329496777;
cosLookup[12882] <= 0.32940625;
cosLookup[12883] <= 0.32931572;
cosLookup[12884] <= 0.329225187;
cosLookup[12885] <= 0.329134651;
cosLookup[12886] <= 0.329044112;
cosLookup[12887] <= 0.32895357;
cosLookup[12888] <= 0.328863025;
cosLookup[12889] <= 0.328772477;
cosLookup[12890] <= 0.328681926;
cosLookup[12891] <= 0.328591371;
cosLookup[12892] <= 0.328500814;
cosLookup[12893] <= 0.328410254;
cosLookup[12894] <= 0.328319691;
cosLookup[12895] <= 0.328229125;
cosLookup[12896] <= 0.328138555;
cosLookup[12897] <= 0.328047983;
cosLookup[12898] <= 0.327957408;
cosLookup[12899] <= 0.32786683;
cosLookup[12900] <= 0.327776248;
cosLookup[12901] <= 0.327685664;
cosLookup[12902] <= 0.327595077;
cosLookup[12903] <= 0.327504486;
cosLookup[12904] <= 0.327413893;
cosLookup[12905] <= 0.327323297;
cosLookup[12906] <= 0.327232697;
cosLookup[12907] <= 0.327142095;
cosLookup[12908] <= 0.327051489;
cosLookup[12909] <= 0.326960881;
cosLookup[12910] <= 0.32687027;
cosLookup[12911] <= 0.326779655;
cosLookup[12912] <= 0.326689038;
cosLookup[12913] <= 0.326598417;
cosLookup[12914] <= 0.326507794;
cosLookup[12915] <= 0.326417168;
cosLookup[12916] <= 0.326326538;
cosLookup[12917] <= 0.326235906;
cosLookup[12918] <= 0.32614527;
cosLookup[12919] <= 0.326054632;
cosLookup[12920] <= 0.32596399;
cosLookup[12921] <= 0.325873346;
cosLookup[12922] <= 0.325782699;
cosLookup[12923] <= 0.325692048;
cosLookup[12924] <= 0.325601395;
cosLookup[12925] <= 0.325510738;
cosLookup[12926] <= 0.325420079;
cosLookup[12927] <= 0.325329417;
cosLookup[12928] <= 0.325238751;
cosLookup[12929] <= 0.325148083;
cosLookup[12930] <= 0.325057412;
cosLookup[12931] <= 0.324966737;
cosLookup[12932] <= 0.32487606;
cosLookup[12933] <= 0.32478538;
cosLookup[12934] <= 0.324694696;
cosLookup[12935] <= 0.32460401;
cosLookup[12936] <= 0.324513321;
cosLookup[12937] <= 0.324422629;
cosLookup[12938] <= 0.324331933;
cosLookup[12939] <= 0.324241235;
cosLookup[12940] <= 0.324150534;
cosLookup[12941] <= 0.32405983;
cosLookup[12942] <= 0.323969123;
cosLookup[12943] <= 0.323878412;
cosLookup[12944] <= 0.323787699;
cosLookup[12945] <= 0.323696983;
cosLookup[12946] <= 0.323606264;
cosLookup[12947] <= 0.323515542;
cosLookup[12948] <= 0.323424817;
cosLookup[12949] <= 0.323334089;
cosLookup[12950] <= 0.323243358;
cosLookup[12951] <= 0.323152624;
cosLookup[12952] <= 0.323061887;
cosLookup[12953] <= 0.322971148;
cosLookup[12954] <= 0.322880405;
cosLookup[12955] <= 0.322789659;
cosLookup[12956] <= 0.32269891;
cosLookup[12957] <= 0.322608158;
cosLookup[12958] <= 0.322517404;
cosLookup[12959] <= 0.322426646;
cosLookup[12960] <= 0.322335885;
cosLookup[12961] <= 0.322245122;
cosLookup[12962] <= 0.322154355;
cosLookup[12963] <= 0.322063586;
cosLookup[12964] <= 0.321972813;
cosLookup[12965] <= 0.321882038;
cosLookup[12966] <= 0.32179126;
cosLookup[12967] <= 0.321700478;
cosLookup[12968] <= 0.321609694;
cosLookup[12969] <= 0.321518907;
cosLookup[12970] <= 0.321428116;
cosLookup[12971] <= 0.321337323;
cosLookup[12972] <= 0.321246527;
cosLookup[12973] <= 0.321155728;
cosLookup[12974] <= 0.321064926;
cosLookup[12975] <= 0.320974121;
cosLookup[12976] <= 0.320883313;
cosLookup[12977] <= 0.320792502;
cosLookup[12978] <= 0.320701688;
cosLookup[12979] <= 0.320610871;
cosLookup[12980] <= 0.320520052;
cosLookup[12981] <= 0.320429229;
cosLookup[12982] <= 0.320338403;
cosLookup[12983] <= 0.320247575;
cosLookup[12984] <= 0.320156743;
cosLookup[12985] <= 0.320065909;
cosLookup[12986] <= 0.319975072;
cosLookup[12987] <= 0.319884231;
cosLookup[12988] <= 0.319793388;
cosLookup[12989] <= 0.319702542;
cosLookup[12990] <= 0.319611693;
cosLookup[12991] <= 0.31952084;
cosLookup[12992] <= 0.319429985;
cosLookup[12993] <= 0.319339127;
cosLookup[12994] <= 0.319248266;
cosLookup[12995] <= 0.319157403;
cosLookup[12996] <= 0.319066536;
cosLookup[12997] <= 0.318975666;
cosLookup[12998] <= 0.318884794;
cosLookup[12999] <= 0.318793918;
cosLookup[13000] <= 0.318703039;
cosLookup[13001] <= 0.318612158;
cosLookup[13002] <= 0.318521274;
cosLookup[13003] <= 0.318430386;
cosLookup[13004] <= 0.318339496;
cosLookup[13005] <= 0.318248603;
cosLookup[13006] <= 0.318157707;
cosLookup[13007] <= 0.318066808;
cosLookup[13008] <= 0.317975906;
cosLookup[13009] <= 0.317885001;
cosLookup[13010] <= 0.317794093;
cosLookup[13011] <= 0.317703183;
cosLookup[13012] <= 0.317612269;
cosLookup[13013] <= 0.317521353;
cosLookup[13014] <= 0.317430433;
cosLookup[13015] <= 0.317339511;
cosLookup[13016] <= 0.317248585;
cosLookup[13017] <= 0.317157657;
cosLookup[13018] <= 0.317066726;
cosLookup[13019] <= 0.316975792;
cosLookup[13020] <= 0.316884855;
cosLookup[13021] <= 0.316793915;
cosLookup[13022] <= 0.316702973;
cosLookup[13023] <= 0.316612027;
cosLookup[13024] <= 0.316521078;
cosLookup[13025] <= 0.316430127;
cosLookup[13026] <= 0.316339172;
cosLookup[13027] <= 0.316248215;
cosLookup[13028] <= 0.316157255;
cosLookup[13029] <= 0.316066292;
cosLookup[13030] <= 0.315975326;
cosLookup[13031] <= 0.315884357;
cosLookup[13032] <= 0.315793385;
cosLookup[13033] <= 0.31570241;
cosLookup[13034] <= 0.315611433;
cosLookup[13035] <= 0.315520452;
cosLookup[13036] <= 0.315429468;
cosLookup[13037] <= 0.315338482;
cosLookup[13038] <= 0.315247493;
cosLookup[13039] <= 0.315156501;
cosLookup[13040] <= 0.315065506;
cosLookup[13041] <= 0.314974508;
cosLookup[13042] <= 0.314883507;
cosLookup[13043] <= 0.314792503;
cosLookup[13044] <= 0.314701497;
cosLookup[13045] <= 0.314610487;
cosLookup[13046] <= 0.314519475;
cosLookup[13047] <= 0.314428459;
cosLookup[13048] <= 0.314337441;
cosLookup[13049] <= 0.31424642;
cosLookup[13050] <= 0.314155396;
cosLookup[13051] <= 0.314064369;
cosLookup[13052] <= 0.313973339;
cosLookup[13053] <= 0.313882307;
cosLookup[13054] <= 0.313791271;
cosLookup[13055] <= 0.313700233;
cosLookup[13056] <= 0.313609192;
cosLookup[13057] <= 0.313518147;
cosLookup[13058] <= 0.3134271;
cosLookup[13059] <= 0.31333605;
cosLookup[13060] <= 0.313244998;
cosLookup[13061] <= 0.313153942;
cosLookup[13062] <= 0.313062883;
cosLookup[13063] <= 0.312971822;
cosLookup[13064] <= 0.312880758;
cosLookup[13065] <= 0.31278969;
cosLookup[13066] <= 0.31269862;
cosLookup[13067] <= 0.312607547;
cosLookup[13068] <= 0.312516472;
cosLookup[13069] <= 0.312425393;
cosLookup[13070] <= 0.312334311;
cosLookup[13071] <= 0.312243227;
cosLookup[13072] <= 0.31215214;
cosLookup[13073] <= 0.312061049;
cosLookup[13074] <= 0.311969956;
cosLookup[13075] <= 0.31187886;
cosLookup[13076] <= 0.311787762;
cosLookup[13077] <= 0.31169666;
cosLookup[13078] <= 0.311605555;
cosLookup[13079] <= 0.311514448;
cosLookup[13080] <= 0.311423338;
cosLookup[13081] <= 0.311332225;
cosLookup[13082] <= 0.311241109;
cosLookup[13083] <= 0.31114999;
cosLookup[13084] <= 0.311058868;
cosLookup[13085] <= 0.310967744;
cosLookup[13086] <= 0.310876616;
cosLookup[13087] <= 0.310785486;
cosLookup[13088] <= 0.310694353;
cosLookup[13089] <= 0.310603217;
cosLookup[13090] <= 0.310512078;
cosLookup[13091] <= 0.310420936;
cosLookup[13092] <= 0.310329792;
cosLookup[13093] <= 0.310238644;
cosLookup[13094] <= 0.310147494;
cosLookup[13095] <= 0.310056341;
cosLookup[13096] <= 0.309965185;
cosLookup[13097] <= 0.309874026;
cosLookup[13098] <= 0.309782865;
cosLookup[13099] <= 0.3096917;
cosLookup[13100] <= 0.309600533;
cosLookup[13101] <= 0.309509363;
cosLookup[13102] <= 0.30941819;
cosLookup[13103] <= 0.309327014;
cosLookup[13104] <= 0.309235835;
cosLookup[13105] <= 0.309144653;
cosLookup[13106] <= 0.309053469;
cosLookup[13107] <= 0.308962282;
cosLookup[13108] <= 0.308871092;
cosLookup[13109] <= 0.308779899;
cosLookup[13110] <= 0.308688703;
cosLookup[13111] <= 0.308597504;
cosLookup[13112] <= 0.308506303;
cosLookup[13113] <= 0.308415099;
cosLookup[13114] <= 0.308323891;
cosLookup[13115] <= 0.308232681;
cosLookup[13116] <= 0.308141469;
cosLookup[13117] <= 0.308050253;
cosLookup[13118] <= 0.307959035;
cosLookup[13119] <= 0.307867813;
cosLookup[13120] <= 0.307776589;
cosLookup[13121] <= 0.307685362;
cosLookup[13122] <= 0.307594133;
cosLookup[13123] <= 0.3075029;
cosLookup[13124] <= 0.307411665;
cosLookup[13125] <= 0.307320426;
cosLookup[13126] <= 0.307229185;
cosLookup[13127] <= 0.307137941;
cosLookup[13128] <= 0.307046695;
cosLookup[13129] <= 0.306955445;
cosLookup[13130] <= 0.306864193;
cosLookup[13131] <= 0.306772938;
cosLookup[13132] <= 0.306681679;
cosLookup[13133] <= 0.306590419;
cosLookup[13134] <= 0.306499155;
cosLookup[13135] <= 0.306407889;
cosLookup[13136] <= 0.306316619;
cosLookup[13137] <= 0.306225347;
cosLookup[13138] <= 0.306134072;
cosLookup[13139] <= 0.306042795;
cosLookup[13140] <= 0.305951514;
cosLookup[13141] <= 0.305860231;
cosLookup[13142] <= 0.305768945;
cosLookup[13143] <= 0.305677656;
cosLookup[13144] <= 0.305586364;
cosLookup[13145] <= 0.305495069;
cosLookup[13146] <= 0.305403772;
cosLookup[13147] <= 0.305312472;
cosLookup[13148] <= 0.305221169;
cosLookup[13149] <= 0.305129863;
cosLookup[13150] <= 0.305038554;
cosLookup[13151] <= 0.304947243;
cosLookup[13152] <= 0.304855928;
cosLookup[13153] <= 0.304764611;
cosLookup[13154] <= 0.304673292;
cosLookup[13155] <= 0.304581969;
cosLookup[13156] <= 0.304490643;
cosLookup[13157] <= 0.304399315;
cosLookup[13158] <= 0.304307984;
cosLookup[13159] <= 0.30421665;
cosLookup[13160] <= 0.304125314;
cosLookup[13161] <= 0.304033974;
cosLookup[13162] <= 0.303942632;
cosLookup[13163] <= 0.303851287;
cosLookup[13164] <= 0.303759939;
cosLookup[13165] <= 0.303668589;
cosLookup[13166] <= 0.303577235;
cosLookup[13167] <= 0.303485879;
cosLookup[13168] <= 0.30339452;
cosLookup[13169] <= 0.303303158;
cosLookup[13170] <= 0.303211794;
cosLookup[13171] <= 0.303120426;
cosLookup[13172] <= 0.303029056;
cosLookup[13173] <= 0.302937683;
cosLookup[13174] <= 0.302846308;
cosLookup[13175] <= 0.302754929;
cosLookup[13176] <= 0.302663548;
cosLookup[13177] <= 0.302572164;
cosLookup[13178] <= 0.302480777;
cosLookup[13179] <= 0.302389388;
cosLookup[13180] <= 0.302297995;
cosLookup[13181] <= 0.3022066;
cosLookup[13182] <= 0.302115202;
cosLookup[13183] <= 0.302023801;
cosLookup[13184] <= 0.301932398;
cosLookup[13185] <= 0.301840992;
cosLookup[13186] <= 0.301749583;
cosLookup[13187] <= 0.301658171;
cosLookup[13188] <= 0.301566756;
cosLookup[13189] <= 0.301475339;
cosLookup[13190] <= 0.301383919;
cosLookup[13191] <= 0.301292496;
cosLookup[13192] <= 0.30120107;
cosLookup[13193] <= 0.301109642;
cosLookup[13194] <= 0.30101821;
cosLookup[13195] <= 0.300926776;
cosLookup[13196] <= 0.30083534;
cosLookup[13197] <= 0.3007439;
cosLookup[13198] <= 0.300652458;
cosLookup[13199] <= 0.300561013;
cosLookup[13200] <= 0.300469565;
cosLookup[13201] <= 0.300378114;
cosLookup[13202] <= 0.300286661;
cosLookup[13203] <= 0.300195205;
cosLookup[13204] <= 0.300103746;
cosLookup[13205] <= 0.300012285;
cosLookup[13206] <= 0.29992082;
cosLookup[13207] <= 0.299829353;
cosLookup[13208] <= 0.299737883;
cosLookup[13209] <= 0.299646411;
cosLookup[13210] <= 0.299554935;
cosLookup[13211] <= 0.299463457;
cosLookup[13212] <= 0.299371976;
cosLookup[13213] <= 0.299280492;
cosLookup[13214] <= 0.299189006;
cosLookup[13215] <= 0.299097517;
cosLookup[13216] <= 0.299006025;
cosLookup[13217] <= 0.29891453;
cosLookup[13218] <= 0.298823033;
cosLookup[13219] <= 0.298731533;
cosLookup[13220] <= 0.29864003;
cosLookup[13221] <= 0.298548524;
cosLookup[13222] <= 0.298457016;
cosLookup[13223] <= 0.298365505;
cosLookup[13224] <= 0.298273991;
cosLookup[13225] <= 0.298182474;
cosLookup[13226] <= 0.298090955;
cosLookup[13227] <= 0.297999433;
cosLookup[13228] <= 0.297907908;
cosLookup[13229] <= 0.29781638;
cosLookup[13230] <= 0.29772485;
cosLookup[13231] <= 0.297633317;
cosLookup[13232] <= 0.297541781;
cosLookup[13233] <= 0.297450243;
cosLookup[13234] <= 0.297358702;
cosLookup[13235] <= 0.297267158;
cosLookup[13236] <= 0.297175611;
cosLookup[13237] <= 0.297084061;
cosLookup[13238] <= 0.296992509;
cosLookup[13239] <= 0.296900954;
cosLookup[13240] <= 0.296809397;
cosLookup[13241] <= 0.296717836;
cosLookup[13242] <= 0.296626273;
cosLookup[13243] <= 0.296534707;
cosLookup[13244] <= 0.296443139;
cosLookup[13245] <= 0.296351568;
cosLookup[13246] <= 0.296259994;
cosLookup[13247] <= 0.296168417;
cosLookup[13248] <= 0.296076837;
cosLookup[13249] <= 0.295985255;
cosLookup[13250] <= 0.29589367;
cosLookup[13251] <= 0.295802083;
cosLookup[13252] <= 0.295710492;
cosLookup[13253] <= 0.295618899;
cosLookup[13254] <= 0.295527304;
cosLookup[13255] <= 0.295435705;
cosLookup[13256] <= 0.295344104;
cosLookup[13257] <= 0.2952525;
cosLookup[13258] <= 0.295160893;
cosLookup[13259] <= 0.295069284;
cosLookup[13260] <= 0.294977672;
cosLookup[13261] <= 0.294886057;
cosLookup[13262] <= 0.29479444;
cosLookup[13263] <= 0.29470282;
cosLookup[13264] <= 0.294611197;
cosLookup[13265] <= 0.294519571;
cosLookup[13266] <= 0.294427943;
cosLookup[13267] <= 0.294336312;
cosLookup[13268] <= 0.294244678;
cosLookup[13269] <= 0.294153042;
cosLookup[13270] <= 0.294061403;
cosLookup[13271] <= 0.293969761;
cosLookup[13272] <= 0.293878116;
cosLookup[13273] <= 0.293786469;
cosLookup[13274] <= 0.293694819;
cosLookup[13275] <= 0.293603166;
cosLookup[13276] <= 0.293511511;
cosLookup[13277] <= 0.293419853;
cosLookup[13278] <= 0.293328192;
cosLookup[13279] <= 0.293236529;
cosLookup[13280] <= 0.293144863;
cosLookup[13281] <= 0.293053194;
cosLookup[13282] <= 0.292961522;
cosLookup[13283] <= 0.292869848;
cosLookup[13284] <= 0.292778171;
cosLookup[13285] <= 0.292686492;
cosLookup[13286] <= 0.29259481;
cosLookup[13287] <= 0.292503125;
cosLookup[13288] <= 0.292411437;
cosLookup[13289] <= 0.292319747;
cosLookup[13290] <= 0.292228053;
cosLookup[13291] <= 0.292136358;
cosLookup[13292] <= 0.292044659;
cosLookup[13293] <= 0.291952958;
cosLookup[13294] <= 0.291861255;
cosLookup[13295] <= 0.291769548;
cosLookup[13296] <= 0.291677839;
cosLookup[13297] <= 0.291586127;
cosLookup[13298] <= 0.291494413;
cosLookup[13299] <= 0.291402695;
cosLookup[13300] <= 0.291310976;
cosLookup[13301] <= 0.291219253;
cosLookup[13302] <= 0.291127528;
cosLookup[13303] <= 0.2910358;
cosLookup[13304] <= 0.290944069;
cosLookup[13305] <= 0.290852336;
cosLookup[13306] <= 0.2907606;
cosLookup[13307] <= 0.290668862;
cosLookup[13308] <= 0.29057712;
cosLookup[13309] <= 0.290485376;
cosLookup[13310] <= 0.29039363;
cosLookup[13311] <= 0.290301881;
cosLookup[13312] <= 0.290210129;
cosLookup[13313] <= 0.290118374;
cosLookup[13314] <= 0.290026617;
cosLookup[13315] <= 0.289934857;
cosLookup[13316] <= 0.289843094;
cosLookup[13317] <= 0.289751329;
cosLookup[13318] <= 0.289659561;
cosLookup[13319] <= 0.28956779;
cosLookup[13320] <= 0.289476017;
cosLookup[13321] <= 0.289384241;
cosLookup[13322] <= 0.289292463;
cosLookup[13323] <= 0.289200681;
cosLookup[13324] <= 0.289108897;
cosLookup[13325] <= 0.289017111;
cosLookup[13326] <= 0.288925322;
cosLookup[13327] <= 0.28883353;
cosLookup[13328] <= 0.288741735;
cosLookup[13329] <= 0.288649938;
cosLookup[13330] <= 0.288558138;
cosLookup[13331] <= 0.288466336;
cosLookup[13332] <= 0.288374531;
cosLookup[13333] <= 0.288282723;
cosLookup[13334] <= 0.288190912;
cosLookup[13335] <= 0.288099099;
cosLookup[13336] <= 0.288007284;
cosLookup[13337] <= 0.287915465;
cosLookup[13338] <= 0.287823644;
cosLookup[13339] <= 0.287731821;
cosLookup[13340] <= 0.287639994;
cosLookup[13341] <= 0.287548165;
cosLookup[13342] <= 0.287456334;
cosLookup[13343] <= 0.287364499;
cosLookup[13344] <= 0.287272663;
cosLookup[13345] <= 0.287180823;
cosLookup[13346] <= 0.287088981;
cosLookup[13347] <= 0.286997136;
cosLookup[13348] <= 0.286905289;
cosLookup[13349] <= 0.286813438;
cosLookup[13350] <= 0.286721586;
cosLookup[13351] <= 0.28662973;
cosLookup[13352] <= 0.286537872;
cosLookup[13353] <= 0.286446012;
cosLookup[13354] <= 0.286354148;
cosLookup[13355] <= 0.286262283;
cosLookup[13356] <= 0.286170414;
cosLookup[13357] <= 0.286078543;
cosLookup[13358] <= 0.285986669;
cosLookup[13359] <= 0.285894793;
cosLookup[13360] <= 0.285802914;
cosLookup[13361] <= 0.285711032;
cosLookup[13362] <= 0.285619148;
cosLookup[13363] <= 0.285527261;
cosLookup[13364] <= 0.285435371;
cosLookup[13365] <= 0.285343479;
cosLookup[13366] <= 0.285251584;
cosLookup[13367] <= 0.285159687;
cosLookup[13368] <= 0.285067787;
cosLookup[13369] <= 0.284975884;
cosLookup[13370] <= 0.284883979;
cosLookup[13371] <= 0.284792071;
cosLookup[13372] <= 0.28470016;
cosLookup[13373] <= 0.284608247;
cosLookup[13374] <= 0.284516332;
cosLookup[13375] <= 0.284424413;
cosLookup[13376] <= 0.284332492;
cosLookup[13377] <= 0.284240569;
cosLookup[13378] <= 0.284148642;
cosLookup[13379] <= 0.284056714;
cosLookup[13380] <= 0.283964782;
cosLookup[13381] <= 0.283872848;
cosLookup[13382] <= 0.283780911;
cosLookup[13383] <= 0.283688972;
cosLookup[13384] <= 0.28359703;
cosLookup[13385] <= 0.283505086;
cosLookup[13386] <= 0.283413139;
cosLookup[13387] <= 0.283321189;
cosLookup[13388] <= 0.283229237;
cosLookup[13389] <= 0.283137282;
cosLookup[13390] <= 0.283045324;
cosLookup[13391] <= 0.282953364;
cosLookup[13392] <= 0.282861402;
cosLookup[13393] <= 0.282769436;
cosLookup[13394] <= 0.282677468;
cosLookup[13395] <= 0.282585498;
cosLookup[13396] <= 0.282493525;
cosLookup[13397] <= 0.282401549;
cosLookup[13398] <= 0.282309571;
cosLookup[13399] <= 0.28221759;
cosLookup[13400] <= 0.282125606;
cosLookup[13401] <= 0.28203362;
cosLookup[13402] <= 0.281941632;
cosLookup[13403] <= 0.28184964;
cosLookup[13404] <= 0.281757647;
cosLookup[13405] <= 0.28166565;
cosLookup[13406] <= 0.281573651;
cosLookup[13407] <= 0.281481649;
cosLookup[13408] <= 0.281389645;
cosLookup[13409] <= 0.281297638;
cosLookup[13410] <= 0.281205629;
cosLookup[13411] <= 0.281113617;
cosLookup[13412] <= 0.281021603;
cosLookup[13413] <= 0.280929585;
cosLookup[13414] <= 0.280837566;
cosLookup[13415] <= 0.280745543;
cosLookup[13416] <= 0.280653519;
cosLookup[13417] <= 0.280561491;
cosLookup[13418] <= 0.280469461;
cosLookup[13419] <= 0.280377428;
cosLookup[13420] <= 0.280285393;
cosLookup[13421] <= 0.280193355;
cosLookup[13422] <= 0.280101315;
cosLookup[13423] <= 0.280009272;
cosLookup[13424] <= 0.279917227;
cosLookup[13425] <= 0.279825179;
cosLookup[13426] <= 0.279733128;
cosLookup[13427] <= 0.279641075;
cosLookup[13428] <= 0.279549019;
cosLookup[13429] <= 0.279456961;
cosLookup[13430] <= 0.2793649;
cosLookup[13431] <= 0.279272836;
cosLookup[13432] <= 0.27918077;
cosLookup[13433] <= 0.279088702;
cosLookup[13434] <= 0.27899663;
cosLookup[13435] <= 0.278904557;
cosLookup[13436] <= 0.27881248;
cosLookup[13437] <= 0.278720401;
cosLookup[13438] <= 0.27862832;
cosLookup[13439] <= 0.278536236;
cosLookup[13440] <= 0.278444149;
cosLookup[13441] <= 0.27835206;
cosLookup[13442] <= 0.278259969;
cosLookup[13443] <= 0.278167874;
cosLookup[13444] <= 0.278075778;
cosLookup[13445] <= 0.277983678;
cosLookup[13446] <= 0.277891576;
cosLookup[13447] <= 0.277799472;
cosLookup[13448] <= 0.277707365;
cosLookup[13449] <= 0.277615255;
cosLookup[13450] <= 0.277523143;
cosLookup[13451] <= 0.277431028;
cosLookup[13452] <= 0.277338911;
cosLookup[13453] <= 0.277246791;
cosLookup[13454] <= 0.277154669;
cosLookup[13455] <= 0.277062544;
cosLookup[13456] <= 0.276970417;
cosLookup[13457] <= 0.276878287;
cosLookup[13458] <= 0.276786154;
cosLookup[13459] <= 0.276694019;
cosLookup[13460] <= 0.276601882;
cosLookup[13461] <= 0.276509742;
cosLookup[13462] <= 0.276417599;
cosLookup[13463] <= 0.276325454;
cosLookup[13464] <= 0.276233306;
cosLookup[13465] <= 0.276141156;
cosLookup[13466] <= 0.276049003;
cosLookup[13467] <= 0.275956847;
cosLookup[13468] <= 0.27586469;
cosLookup[13469] <= 0.275772529;
cosLookup[13470] <= 0.275680366;
cosLookup[13471] <= 0.275588201;
cosLookup[13472] <= 0.275496033;
cosLookup[13473] <= 0.275403862;
cosLookup[13474] <= 0.275311689;
cosLookup[13475] <= 0.275219513;
cosLookup[13476] <= 0.275127335;
cosLookup[13477] <= 0.275035154;
cosLookup[13478] <= 0.274942971;
cosLookup[13479] <= 0.274850785;
cosLookup[13480] <= 0.274758597;
cosLookup[13481] <= 0.274666406;
cosLookup[13482] <= 0.274574213;
cosLookup[13483] <= 0.274482017;
cosLookup[13484] <= 0.274389819;
cosLookup[13485] <= 0.274297618;
cosLookup[13486] <= 0.274205414;
cosLookup[13487] <= 0.274113208;
cosLookup[13488] <= 0.274021;
cosLookup[13489] <= 0.273928789;
cosLookup[13490] <= 0.273836575;
cosLookup[13491] <= 0.273744359;
cosLookup[13492] <= 0.273652141;
cosLookup[13493] <= 0.27355992;
cosLookup[13494] <= 0.273467696;
cosLookup[13495] <= 0.27337547;
cosLookup[13496] <= 0.273283241;
cosLookup[13497] <= 0.27319101;
cosLookup[13498] <= 0.273098777;
cosLookup[13499] <= 0.27300654;
cosLookup[13500] <= 0.272914302;
cosLookup[13501] <= 0.272822061;
cosLookup[13502] <= 0.272729817;
cosLookup[13503] <= 0.272637571;
cosLookup[13504] <= 0.272545322;
cosLookup[13505] <= 0.272453071;
cosLookup[13506] <= 0.272360817;
cosLookup[13507] <= 0.272268561;
cosLookup[13508] <= 0.272176302;
cosLookup[13509] <= 0.272084041;
cosLookup[13510] <= 0.271991778;
cosLookup[13511] <= 0.271899511;
cosLookup[13512] <= 0.271807243;
cosLookup[13513] <= 0.271714971;
cosLookup[13514] <= 0.271622698;
cosLookup[13515] <= 0.271530422;
cosLookup[13516] <= 0.271438143;
cosLookup[13517] <= 0.271345862;
cosLookup[13518] <= 0.271253578;
cosLookup[13519] <= 0.271161292;
cosLookup[13520] <= 0.271069003;
cosLookup[13521] <= 0.270976712;
cosLookup[13522] <= 0.270884418;
cosLookup[13523] <= 0.270792122;
cosLookup[13524] <= 0.270699824;
cosLookup[13525] <= 0.270607522;
cosLookup[13526] <= 0.270515219;
cosLookup[13527] <= 0.270422913;
cosLookup[13528] <= 0.270330604;
cosLookup[13529] <= 0.270238293;
cosLookup[13530] <= 0.27014598;
cosLookup[13531] <= 0.270053664;
cosLookup[13532] <= 0.269961345;
cosLookup[13533] <= 0.269869024;
cosLookup[13534] <= 0.269776701;
cosLookup[13535] <= 0.269684375;
cosLookup[13536] <= 0.269592046;
cosLookup[13537] <= 0.269499715;
cosLookup[13538] <= 0.269407382;
cosLookup[13539] <= 0.269315046;
cosLookup[13540] <= 0.269222708;
cosLookup[13541] <= 0.269130367;
cosLookup[13542] <= 0.269038024;
cosLookup[13543] <= 0.268945678;
cosLookup[13544] <= 0.26885333;
cosLookup[13545] <= 0.268760979;
cosLookup[13546] <= 0.268668626;
cosLookup[13547] <= 0.26857627;
cosLookup[13548] <= 0.268483912;
cosLookup[13549] <= 0.268391551;
cosLookup[13550] <= 0.268299188;
cosLookup[13551] <= 0.268206823;
cosLookup[13552] <= 0.268114455;
cosLookup[13553] <= 0.268022084;
cosLookup[13554] <= 0.267929711;
cosLookup[13555] <= 0.267837336;
cosLookup[13556] <= 0.267744958;
cosLookup[13557] <= 0.267652578;
cosLookup[13558] <= 0.267560195;
cosLookup[13559] <= 0.26746781;
cosLookup[13560] <= 0.267375422;
cosLookup[13561] <= 0.267283032;
cosLookup[13562] <= 0.26719064;
cosLookup[13563] <= 0.267098245;
cosLookup[13564] <= 0.267005847;
cosLookup[13565] <= 0.266913447;
cosLookup[13566] <= 0.266821045;
cosLookup[13567] <= 0.26672864;
cosLookup[13568] <= 0.266636232;
cosLookup[13569] <= 0.266543823;
cosLookup[13570] <= 0.266451411;
cosLookup[13571] <= 0.266358996;
cosLookup[13572] <= 0.266266579;
cosLookup[13573] <= 0.266174159;
cosLookup[13574] <= 0.266081737;
cosLookup[13575] <= 0.265989313;
cosLookup[13576] <= 0.265896886;
cosLookup[13577] <= 0.265804456;
cosLookup[13578] <= 0.265712025;
cosLookup[13579] <= 0.26561959;
cosLookup[13580] <= 0.265527154;
cosLookup[13581] <= 0.265434715;
cosLookup[13582] <= 0.265342273;
cosLookup[13583] <= 0.265249829;
cosLookup[13584] <= 0.265157383;
cosLookup[13585] <= 0.265064934;
cosLookup[13586] <= 0.264972482;
cosLookup[13587] <= 0.264880029;
cosLookup[13588] <= 0.264787573;
cosLookup[13589] <= 0.264695114;
cosLookup[13590] <= 0.264602653;
cosLookup[13591] <= 0.264510189;
cosLookup[13592] <= 0.264417723;
cosLookup[13593] <= 0.264325255;
cosLookup[13594] <= 0.264232784;
cosLookup[13595] <= 0.264140311;
cosLookup[13596] <= 0.264047836;
cosLookup[13597] <= 0.263955357;
cosLookup[13598] <= 0.263862877;
cosLookup[13599] <= 0.263770394;
cosLookup[13600] <= 0.263677909;
cosLookup[13601] <= 0.263585421;
cosLookup[13602] <= 0.263492931;
cosLookup[13603] <= 0.263400438;
cosLookup[13604] <= 0.263307943;
cosLookup[13605] <= 0.263215446;
cosLookup[13606] <= 0.263122946;
cosLookup[13607] <= 0.263030444;
cosLookup[13608] <= 0.262937939;
cosLookup[13609] <= 0.262845432;
cosLookup[13610] <= 0.262752922;
cosLookup[13611] <= 0.26266041;
cosLookup[13612] <= 0.262567896;
cosLookup[13613] <= 0.262475379;
cosLookup[13614] <= 0.26238286;
cosLookup[13615] <= 0.262290338;
cosLookup[13616] <= 0.262197814;
cosLookup[13617] <= 0.262105288;
cosLookup[13618] <= 0.262012759;
cosLookup[13619] <= 0.261920228;
cosLookup[13620] <= 0.261827694;
cosLookup[13621] <= 0.261735158;
cosLookup[13622] <= 0.26164262;
cosLookup[13623] <= 0.261550079;
cosLookup[13624] <= 0.261457536;
cosLookup[13625] <= 0.26136499;
cosLookup[13626] <= 0.261272442;
cosLookup[13627] <= 0.261179891;
cosLookup[13628] <= 0.261087338;
cosLookup[13629] <= 0.260994783;
cosLookup[13630] <= 0.260902225;
cosLookup[13631] <= 0.260809665;
cosLookup[13632] <= 0.260717103;
cosLookup[13633] <= 0.260624538;
cosLookup[13634] <= 0.260531971;
cosLookup[13635] <= 0.260439401;
cosLookup[13636] <= 0.260346829;
cosLookup[13637] <= 0.260254255;
cosLookup[13638] <= 0.260161678;
cosLookup[13639] <= 0.260069098;
cosLookup[13640] <= 0.259976517;
cosLookup[13641] <= 0.259883933;
cosLookup[13642] <= 0.259791346;
cosLookup[13643] <= 0.259698758;
cosLookup[13644] <= 0.259606166;
cosLookup[13645] <= 0.259513573;
cosLookup[13646] <= 0.259420977;
cosLookup[13647] <= 0.259328379;
cosLookup[13648] <= 0.259235778;
cosLookup[13649] <= 0.259143175;
cosLookup[13650] <= 0.259050569;
cosLookup[13651] <= 0.258957961;
cosLookup[13652] <= 0.258865351;
cosLookup[13653] <= 0.258772738;
cosLookup[13654] <= 0.258680123;
cosLookup[13655] <= 0.258587506;
cosLookup[13656] <= 0.258494886;
cosLookup[13657] <= 0.258402264;
cosLookup[13658] <= 0.25830964;
cosLookup[13659] <= 0.258217013;
cosLookup[13660] <= 0.258124384;
cosLookup[13661] <= 0.258031752;
cosLookup[13662] <= 0.257939118;
cosLookup[13663] <= 0.257846481;
cosLookup[13664] <= 0.257753843;
cosLookup[13665] <= 0.257661202;
cosLookup[13666] <= 0.257568558;
cosLookup[13667] <= 0.257475912;
cosLookup[13668] <= 0.257383264;
cosLookup[13669] <= 0.257290613;
cosLookup[13670] <= 0.25719796;
cosLookup[13671] <= 0.257105305;
cosLookup[13672] <= 0.257012647;
cosLookup[13673] <= 0.256919987;
cosLookup[13674] <= 0.256827325;
cosLookup[13675] <= 0.25673466;
cosLookup[13676] <= 0.256641993;
cosLookup[13677] <= 0.256549324;
cosLookup[13678] <= 0.256456652;
cosLookup[13679] <= 0.256363978;
cosLookup[13680] <= 0.256271301;
cosLookup[13681] <= 0.256178622;
cosLookup[13682] <= 0.256085941;
cosLookup[13683] <= 0.255993257;
cosLookup[13684] <= 0.255900571;
cosLookup[13685] <= 0.255807883;
cosLookup[13686] <= 0.255715192;
cosLookup[13687] <= 0.255622499;
cosLookup[13688] <= 0.255529804;
cosLookup[13689] <= 0.255437106;
cosLookup[13690] <= 0.255344406;
cosLookup[13691] <= 0.255251704;
cosLookup[13692] <= 0.255158999;
cosLookup[13693] <= 0.255066292;
cosLookup[13694] <= 0.254973582;
cosLookup[13695] <= 0.25488087;
cosLookup[13696] <= 0.254788156;
cosLookup[13697] <= 0.25469544;
cosLookup[13698] <= 0.254602721;
cosLookup[13699] <= 0.25451;
cosLookup[13700] <= 0.254417276;
cosLookup[13701] <= 0.25432455;
cosLookup[13702] <= 0.254231822;
cosLookup[13703] <= 0.254139092;
cosLookup[13704] <= 0.254046359;
cosLookup[13705] <= 0.253953624;
cosLookup[13706] <= 0.253860886;
cosLookup[13707] <= 0.253768146;
cosLookup[13708] <= 0.253675404;
cosLookup[13709] <= 0.253582659;
cosLookup[13710] <= 0.253489913;
cosLookup[13711] <= 0.253397163;
cosLookup[13712] <= 0.253304412;
cosLookup[13713] <= 0.253211658;
cosLookup[13714] <= 0.253118902;
cosLookup[13715] <= 0.253026143;
cosLookup[13716] <= 0.252933382;
cosLookup[13717] <= 0.252840619;
cosLookup[13718] <= 0.252747854;
cosLookup[13719] <= 0.252655086;
cosLookup[13720] <= 0.252562316;
cosLookup[13721] <= 0.252469543;
cosLookup[13722] <= 0.252376769;
cosLookup[13723] <= 0.252283991;
cosLookup[13724] <= 0.252191212;
cosLookup[13725] <= 0.25209843;
cosLookup[13726] <= 0.252005646;
cosLookup[13727] <= 0.25191286;
cosLookup[13728] <= 0.251820071;
cosLookup[13729] <= 0.25172728;
cosLookup[13730] <= 0.251634487;
cosLookup[13731] <= 0.251541691;
cosLookup[13732] <= 0.251448893;
cosLookup[13733] <= 0.251356093;
cosLookup[13734] <= 0.251263291;
cosLookup[13735] <= 0.251170486;
cosLookup[13736] <= 0.251077679;
cosLookup[13737] <= 0.250984869;
cosLookup[13738] <= 0.250892057;
cosLookup[13739] <= 0.250799243;
cosLookup[13740] <= 0.250706427;
cosLookup[13741] <= 0.250613608;
cosLookup[13742] <= 0.250520787;
cosLookup[13743] <= 0.250427964;
cosLookup[13744] <= 0.250335138;
cosLookup[13745] <= 0.25024231;
cosLookup[13746] <= 0.25014948;
cosLookup[13747] <= 0.250056647;
cosLookup[13748] <= 0.249963813;
cosLookup[13749] <= 0.249870975;
cosLookup[13750] <= 0.249778136;
cosLookup[13751] <= 0.249685294;
cosLookup[13752] <= 0.24959245;
cosLookup[13753] <= 0.249499604;
cosLookup[13754] <= 0.249406755;
cosLookup[13755] <= 0.249313905;
cosLookup[13756] <= 0.249221051;
cosLookup[13757] <= 0.249128196;
cosLookup[13758] <= 0.249035338;
cosLookup[13759] <= 0.248942478;
cosLookup[13760] <= 0.248849616;
cosLookup[13761] <= 0.248756751;
cosLookup[13762] <= 0.248663884;
cosLookup[13763] <= 0.248571015;
cosLookup[13764] <= 0.248478144;
cosLookup[13765] <= 0.24838527;
cosLookup[13766] <= 0.248292394;
cosLookup[13767] <= 0.248199515;
cosLookup[13768] <= 0.248106635;
cosLookup[13769] <= 0.248013752;
cosLookup[13770] <= 0.247920867;
cosLookup[13771] <= 0.247827979;
cosLookup[13772] <= 0.247735089;
cosLookup[13773] <= 0.247642197;
cosLookup[13774] <= 0.247549303;
cosLookup[13775] <= 0.247456407;
cosLookup[13776] <= 0.247363508;
cosLookup[13777] <= 0.247270607;
cosLookup[13778] <= 0.247177703;
cosLookup[13779] <= 0.247084798;
cosLookup[13780] <= 0.24699189;
cosLookup[13781] <= 0.24689898;
cosLookup[13782] <= 0.246806067;
cosLookup[13783] <= 0.246713152;
cosLookup[13784] <= 0.246620235;
cosLookup[13785] <= 0.246527316;
cosLookup[13786] <= 0.246434394;
cosLookup[13787] <= 0.246341471;
cosLookup[13788] <= 0.246248545;
cosLookup[13789] <= 0.246155616;
cosLookup[13790] <= 0.246062686;
cosLookup[13791] <= 0.245969753;
cosLookup[13792] <= 0.245876818;
cosLookup[13793] <= 0.24578388;
cosLookup[13794] <= 0.245690941;
cosLookup[13795] <= 0.245597999;
cosLookup[13796] <= 0.245505055;
cosLookup[13797] <= 0.245412108;
cosLookup[13798] <= 0.24531916;
cosLookup[13799] <= 0.245226209;
cosLookup[13800] <= 0.245133255;
cosLookup[13801] <= 0.2450403;
cosLookup[13802] <= 0.244947342;
cosLookup[13803] <= 0.244854382;
cosLookup[13804] <= 0.24476142;
cosLookup[13805] <= 0.244668456;
cosLookup[13806] <= 0.244575489;
cosLookup[13807] <= 0.24448252;
cosLookup[13808] <= 0.244389549;
cosLookup[13809] <= 0.244296576;
cosLookup[13810] <= 0.2442036;
cosLookup[13811] <= 0.244110622;
cosLookup[13812] <= 0.244017642;
cosLookup[13813] <= 0.243924659;
cosLookup[13814] <= 0.243831675;
cosLookup[13815] <= 0.243738688;
cosLookup[13816] <= 0.243645699;
cosLookup[13817] <= 0.243552707;
cosLookup[13818] <= 0.243459714;
cosLookup[13819] <= 0.243366718;
cosLookup[13820] <= 0.24327372;
cosLookup[13821] <= 0.243180719;
cosLookup[13822] <= 0.243087717;
cosLookup[13823] <= 0.242994712;
cosLookup[13824] <= 0.242901705;
cosLookup[13825] <= 0.242808696;
cosLookup[13826] <= 0.242715684;
cosLookup[13827] <= 0.242622671;
cosLookup[13828] <= 0.242529655;
cosLookup[13829] <= 0.242436636;
cosLookup[13830] <= 0.242343616;
cosLookup[13831] <= 0.242250593;
cosLookup[13832] <= 0.242157569;
cosLookup[13833] <= 0.242064541;
cosLookup[13834] <= 0.241971512;
cosLookup[13835] <= 0.241878481;
cosLookup[13836] <= 0.241785447;
cosLookup[13837] <= 0.241692411;
cosLookup[13838] <= 0.241599373;
cosLookup[13839] <= 0.241506332;
cosLookup[13840] <= 0.24141329;
cosLookup[13841] <= 0.241320245;
cosLookup[13842] <= 0.241227198;
cosLookup[13843] <= 0.241134148;
cosLookup[13844] <= 0.241041097;
cosLookup[13845] <= 0.240948043;
cosLookup[13846] <= 0.240854987;
cosLookup[13847] <= 0.240761929;
cosLookup[13848] <= 0.240668869;
cosLookup[13849] <= 0.240575806;
cosLookup[13850] <= 0.240482741;
cosLookup[13851] <= 0.240389674;
cosLookup[13852] <= 0.240296605;
cosLookup[13853] <= 0.240203533;
cosLookup[13854] <= 0.24011046;
cosLookup[13855] <= 0.240017384;
cosLookup[13856] <= 0.239924306;
cosLookup[13857] <= 0.239831226;
cosLookup[13858] <= 0.239738143;
cosLookup[13859] <= 0.239645059;
cosLookup[13860] <= 0.239551972;
cosLookup[13861] <= 0.239458883;
cosLookup[13862] <= 0.239365791;
cosLookup[13863] <= 0.239272698;
cosLookup[13864] <= 0.239179602;
cosLookup[13865] <= 0.239086504;
cosLookup[13866] <= 0.238993404;
cosLookup[13867] <= 0.238900302;
cosLookup[13868] <= 0.238807197;
cosLookup[13869] <= 0.238714091;
cosLookup[13870] <= 0.238620982;
cosLookup[13871] <= 0.238527871;
cosLookup[13872] <= 0.238434758;
cosLookup[13873] <= 0.238341642;
cosLookup[13874] <= 0.238248525;
cosLookup[13875] <= 0.238155405;
cosLookup[13876] <= 0.238062283;
cosLookup[13877] <= 0.237969159;
cosLookup[13878] <= 0.237876032;
cosLookup[13879] <= 0.237782904;
cosLookup[13880] <= 0.237689773;
cosLookup[13881] <= 0.23759664;
cosLookup[13882] <= 0.237503505;
cosLookup[13883] <= 0.237410367;
cosLookup[13884] <= 0.237317228;
cosLookup[13885] <= 0.237224086;
cosLookup[13886] <= 0.237130942;
cosLookup[13887] <= 0.237037796;
cosLookup[13888] <= 0.236944648;
cosLookup[13889] <= 0.236851498;
cosLookup[13890] <= 0.236758345;
cosLookup[13891] <= 0.23666519;
cosLookup[13892] <= 0.236572034;
cosLookup[13893] <= 0.236478874;
cosLookup[13894] <= 0.236385713;
cosLookup[13895] <= 0.23629255;
cosLookup[13896] <= 0.236199384;
cosLookup[13897] <= 0.236106216;
cosLookup[13898] <= 0.236013046;
cosLookup[13899] <= 0.235919874;
cosLookup[13900] <= 0.2358267;
cosLookup[13901] <= 0.235733524;
cosLookup[13902] <= 0.235640345;
cosLookup[13903] <= 0.235547164;
cosLookup[13904] <= 0.235453981;
cosLookup[13905] <= 0.235360796;
cosLookup[13906] <= 0.235267609;
cosLookup[13907] <= 0.235174419;
cosLookup[13908] <= 0.235081228;
cosLookup[13909] <= 0.234988034;
cosLookup[13910] <= 0.234894838;
cosLookup[13911] <= 0.23480164;
cosLookup[13912] <= 0.23470844;
cosLookup[13913] <= 0.234615237;
cosLookup[13914] <= 0.234522033;
cosLookup[13915] <= 0.234428826;
cosLookup[13916] <= 0.234335617;
cosLookup[13917] <= 0.234242406;
cosLookup[13918] <= 0.234149193;
cosLookup[13919] <= 0.234055977;
cosLookup[13920] <= 0.23396276;
cosLookup[13921] <= 0.23386954;
cosLookup[13922] <= 0.233776319;
cosLookup[13923] <= 0.233683095;
cosLookup[13924] <= 0.233589869;
cosLookup[13925] <= 0.23349664;
cosLookup[13926] <= 0.23340341;
cosLookup[13927] <= 0.233310177;
cosLookup[13928] <= 0.233216943;
cosLookup[13929] <= 0.233123706;
cosLookup[13930] <= 0.233030467;
cosLookup[13931] <= 0.232937226;
cosLookup[13932] <= 0.232843983;
cosLookup[13933] <= 0.232750737;
cosLookup[13934] <= 0.23265749;
cosLookup[13935] <= 0.23256424;
cosLookup[13936] <= 0.232470988;
cosLookup[13937] <= 0.232377734;
cosLookup[13938] <= 0.232284478;
cosLookup[13939] <= 0.23219122;
cosLookup[13940] <= 0.23209796;
cosLookup[13941] <= 0.232004697;
cosLookup[13942] <= 0.231911433;
cosLookup[13943] <= 0.231818166;
cosLookup[13944] <= 0.231724897;
cosLookup[13945] <= 0.231631626;
cosLookup[13946] <= 0.231538353;
cosLookup[13947] <= 0.231445078;
cosLookup[13948] <= 0.2313518;
cosLookup[13949] <= 0.231258521;
cosLookup[13950] <= 0.231165239;
cosLookup[13951] <= 0.231071955;
cosLookup[13952] <= 0.230978669;
cosLookup[13953] <= 0.230885381;
cosLookup[13954] <= 0.230792091;
cosLookup[13955] <= 0.230698799;
cosLookup[13956] <= 0.230605505;
cosLookup[13957] <= 0.230512208;
cosLookup[13958] <= 0.230418909;
cosLookup[13959] <= 0.230325609;
cosLookup[13960] <= 0.230232306;
cosLookup[13961] <= 0.230139001;
cosLookup[13962] <= 0.230045694;
cosLookup[13963] <= 0.229952385;
cosLookup[13964] <= 0.229859073;
cosLookup[13965] <= 0.22976576;
cosLookup[13966] <= 0.229672444;
cosLookup[13967] <= 0.229579127;
cosLookup[13968] <= 0.229485807;
cosLookup[13969] <= 0.229392485;
cosLookup[13970] <= 0.229299161;
cosLookup[13971] <= 0.229205835;
cosLookup[13972] <= 0.229112507;
cosLookup[13973] <= 0.229019177;
cosLookup[13974] <= 0.228925844;
cosLookup[13975] <= 0.22883251;
cosLookup[13976] <= 0.228739173;
cosLookup[13977] <= 0.228645834;
cosLookup[13978] <= 0.228552493;
cosLookup[13979] <= 0.228459151;
cosLookup[13980] <= 0.228365806;
cosLookup[13981] <= 0.228272458;
cosLookup[13982] <= 0.228179109;
cosLookup[13983] <= 0.228085758;
cosLookup[13984] <= 0.227992404;
cosLookup[13985] <= 0.227899049;
cosLookup[13986] <= 0.227805691;
cosLookup[13987] <= 0.227712332;
cosLookup[13988] <= 0.22761897;
cosLookup[13989] <= 0.227525606;
cosLookup[13990] <= 0.22743224;
cosLookup[13991] <= 0.227338872;
cosLookup[13992] <= 0.227245502;
cosLookup[13993] <= 0.22715213;
cosLookup[13994] <= 0.227058755;
cosLookup[13995] <= 0.226965379;
cosLookup[13996] <= 0.226872;
cosLookup[13997] <= 0.22677862;
cosLookup[13998] <= 0.226685237;
cosLookup[13999] <= 0.226591852;
cosLookup[14000] <= 0.226498465;
cosLookup[14001] <= 0.226405076;
cosLookup[14002] <= 0.226311685;
cosLookup[14003] <= 0.226218292;
cosLookup[14004] <= 0.226124897;
cosLookup[14005] <= 0.2260315;
cosLookup[14006] <= 0.225938101;
cosLookup[14007] <= 0.225844699;
cosLookup[14008] <= 0.225751296;
cosLookup[14009] <= 0.22565789;
cosLookup[14010] <= 0.225564483;
cosLookup[14011] <= 0.225471073;
cosLookup[14012] <= 0.225377661;
cosLookup[14013] <= 0.225284247;
cosLookup[14014] <= 0.225190831;
cosLookup[14015] <= 0.225097413;
cosLookup[14016] <= 0.225003993;
cosLookup[14017] <= 0.224910571;
cosLookup[14018] <= 0.224817147;
cosLookup[14019] <= 0.224723721;
cosLookup[14020] <= 0.224630292;
cosLookup[14021] <= 0.224536862;
cosLookup[14022] <= 0.22444343;
cosLookup[14023] <= 0.224349995;
cosLookup[14024] <= 0.224256558;
cosLookup[14025] <= 0.22416312;
cosLookup[14026] <= 0.224069679;
cosLookup[14027] <= 0.223976236;
cosLookup[14028] <= 0.223882792;
cosLookup[14029] <= 0.223789345;
cosLookup[14030] <= 0.223695896;
cosLookup[14031] <= 0.223602445;
cosLookup[14032] <= 0.223508992;
cosLookup[14033] <= 0.223415537;
cosLookup[14034] <= 0.223322079;
cosLookup[14035] <= 0.22322862;
cosLookup[14036] <= 0.223135159;
cosLookup[14037] <= 0.223041696;
cosLookup[14038] <= 0.22294823;
cosLookup[14039] <= 0.222854763;
cosLookup[14040] <= 0.222761293;
cosLookup[14041] <= 0.222667822;
cosLookup[14042] <= 0.222574348;
cosLookup[14043] <= 0.222480873;
cosLookup[14044] <= 0.222387395;
cosLookup[14045] <= 0.222293915;
cosLookup[14046] <= 0.222200434;
cosLookup[14047] <= 0.22210695;
cosLookup[14048] <= 0.222013464;
cosLookup[14049] <= 0.221919976;
cosLookup[14050] <= 0.221826486;
cosLookup[14051] <= 0.221732994;
cosLookup[14052] <= 0.2216395;
cosLookup[14053] <= 0.221546004;
cosLookup[14054] <= 0.221452506;
cosLookup[14055] <= 0.221359006;
cosLookup[14056] <= 0.221265504;
cosLookup[14057] <= 0.221172;
cosLookup[14058] <= 0.221078494;
cosLookup[14059] <= 0.220984986;
cosLookup[14060] <= 0.220891475;
cosLookup[14061] <= 0.220797963;
cosLookup[14062] <= 0.220704449;
cosLookup[14063] <= 0.220610932;
cosLookup[14064] <= 0.220517414;
cosLookup[14065] <= 0.220423894;
cosLookup[14066] <= 0.220330371;
cosLookup[14067] <= 0.220236847;
cosLookup[14068] <= 0.22014332;
cosLookup[14069] <= 0.220049792;
cosLookup[14070] <= 0.219956261;
cosLookup[14071] <= 0.219862729;
cosLookup[14072] <= 0.219769194;
cosLookup[14073] <= 0.219675657;
cosLookup[14074] <= 0.219582119;
cosLookup[14075] <= 0.219488578;
cosLookup[14076] <= 0.219395036;
cosLookup[14077] <= 0.219301491;
cosLookup[14078] <= 0.219207944;
cosLookup[14079] <= 0.219114396;
cosLookup[14080] <= 0.219020845;
cosLookup[14081] <= 0.218927292;
cosLookup[14082] <= 0.218833737;
cosLookup[14083] <= 0.218740181;
cosLookup[14084] <= 0.218646622;
cosLookup[14085] <= 0.218553061;
cosLookup[14086] <= 0.218459498;
cosLookup[14087] <= 0.218365934;
cosLookup[14088] <= 0.218272367;
cosLookup[14089] <= 0.218178798;
cosLookup[14090] <= 0.218085227;
cosLookup[14091] <= 0.217991654;
cosLookup[14092] <= 0.21789808;
cosLookup[14093] <= 0.217804503;
cosLookup[14094] <= 0.217710924;
cosLookup[14095] <= 0.217617343;
cosLookup[14096] <= 0.21752376;
cosLookup[14097] <= 0.217430176;
cosLookup[14098] <= 0.217336589;
cosLookup[14099] <= 0.217243;
cosLookup[14100] <= 0.217149409;
cosLookup[14101] <= 0.217055816;
cosLookup[14102] <= 0.216962222;
cosLookup[14103] <= 0.216868625;
cosLookup[14104] <= 0.216775026;
cosLookup[14105] <= 0.216681425;
cosLookup[14106] <= 0.216587822;
cosLookup[14107] <= 0.216494218;
cosLookup[14108] <= 0.216400611;
cosLookup[14109] <= 0.216307002;
cosLookup[14110] <= 0.216213391;
cosLookup[14111] <= 0.216119779;
cosLookup[14112] <= 0.216026164;
cosLookup[14113] <= 0.215932547;
cosLookup[14114] <= 0.215838929;
cosLookup[14115] <= 0.215745308;
cosLookup[14116] <= 0.215651685;
cosLookup[14117] <= 0.215558061;
cosLookup[14118] <= 0.215464434;
cosLookup[14119] <= 0.215370805;
cosLookup[14120] <= 0.215277175;
cosLookup[14121] <= 0.215183542;
cosLookup[14122] <= 0.215089908;
cosLookup[14123] <= 0.214996271;
cosLookup[14124] <= 0.214902633;
cosLookup[14125] <= 0.214808992;
cosLookup[14126] <= 0.21471535;
cosLookup[14127] <= 0.214621706;
cosLookup[14128] <= 0.214528059;
cosLookup[14129] <= 0.214434411;
cosLookup[14130] <= 0.21434076;
cosLookup[14131] <= 0.214247108;
cosLookup[14132] <= 0.214153454;
cosLookup[14133] <= 0.214059798;
cosLookup[14134] <= 0.21396614;
cosLookup[14135] <= 0.213872479;
cosLookup[14136] <= 0.213778817;
cosLookup[14137] <= 0.213685153;
cosLookup[14138] <= 0.213591487;
cosLookup[14139] <= 0.213497819;
cosLookup[14140] <= 0.213404149;
cosLookup[14141] <= 0.213310477;
cosLookup[14142] <= 0.213216803;
cosLookup[14143] <= 0.213123127;
cosLookup[14144] <= 0.213029449;
cosLookup[14145] <= 0.21293577;
cosLookup[14146] <= 0.212842088;
cosLookup[14147] <= 0.212748404;
cosLookup[14148] <= 0.212654719;
cosLookup[14149] <= 0.212561031;
cosLookup[14150] <= 0.212467341;
cosLookup[14151] <= 0.21237365;
cosLookup[14152] <= 0.212279956;
cosLookup[14153] <= 0.212186261;
cosLookup[14154] <= 0.212092564;
cosLookup[14155] <= 0.211998864;
cosLookup[14156] <= 0.211905163;
cosLookup[14157] <= 0.21181146;
cosLookup[14158] <= 0.211717755;
cosLookup[14159] <= 0.211624048;
cosLookup[14160] <= 0.211530338;
cosLookup[14161] <= 0.211436627;
cosLookup[14162] <= 0.211342915;
cosLookup[14163] <= 0.2112492;
cosLookup[14164] <= 0.211155483;
cosLookup[14165] <= 0.211061764;
cosLookup[14166] <= 0.210968043;
cosLookup[14167] <= 0.210874321;
cosLookup[14168] <= 0.210780596;
cosLookup[14169] <= 0.21068687;
cosLookup[14170] <= 0.210593141;
cosLookup[14171] <= 0.210499411;
cosLookup[14172] <= 0.210405678;
cosLookup[14173] <= 0.210311944;
cosLookup[14174] <= 0.210218208;
cosLookup[14175] <= 0.21012447;
cosLookup[14176] <= 0.21003073;
cosLookup[14177] <= 0.209936988;
cosLookup[14178] <= 0.209843244;
cosLookup[14179] <= 0.209749498;
cosLookup[14180] <= 0.20965575;
cosLookup[14181] <= 0.209562;
cosLookup[14182] <= 0.209468249;
cosLookup[14183] <= 0.209374495;
cosLookup[14184] <= 0.20928074;
cosLookup[14185] <= 0.209186982;
cosLookup[14186] <= 0.209093223;
cosLookup[14187] <= 0.208999462;
cosLookup[14188] <= 0.208905698;
cosLookup[14189] <= 0.208811933;
cosLookup[14190] <= 0.208718166;
cosLookup[14191] <= 0.208624397;
cosLookup[14192] <= 0.208530627;
cosLookup[14193] <= 0.208436854;
cosLookup[14194] <= 0.208343079;
cosLookup[14195] <= 0.208249302;
cosLookup[14196] <= 0.208155524;
cosLookup[14197] <= 0.208061743;
cosLookup[14198] <= 0.207967961;
cosLookup[14199] <= 0.207874177;
cosLookup[14200] <= 0.207780391;
cosLookup[14201] <= 0.207686603;
cosLookup[14202] <= 0.207592813;
cosLookup[14203] <= 0.207499021;
cosLookup[14204] <= 0.207405227;
cosLookup[14205] <= 0.207311431;
cosLookup[14206] <= 0.207217634;
cosLookup[14207] <= 0.207123834;
cosLookup[14208] <= 0.207030033;
cosLookup[14209] <= 0.206936229;
cosLookup[14210] <= 0.206842424;
cosLookup[14211] <= 0.206748617;
cosLookup[14212] <= 0.206654808;
cosLookup[14213] <= 0.206560997;
cosLookup[14214] <= 0.206467184;
cosLookup[14215] <= 0.206373369;
cosLookup[14216] <= 0.206279553;
cosLookup[14217] <= 0.206185734;
cosLookup[14218] <= 0.206091914;
cosLookup[14219] <= 0.205998092;
cosLookup[14220] <= 0.205904267;
cosLookup[14221] <= 0.205810441;
cosLookup[14222] <= 0.205716613;
cosLookup[14223] <= 0.205622783;
cosLookup[14224] <= 0.205528952;
cosLookup[14225] <= 0.205435118;
cosLookup[14226] <= 0.205341282;
cosLookup[14227] <= 0.205247445;
cosLookup[14228] <= 0.205153606;
cosLookup[14229] <= 0.205059764;
cosLookup[14230] <= 0.204965921;
cosLookup[14231] <= 0.204872076;
cosLookup[14232] <= 0.204778229;
cosLookup[14233] <= 0.204684381;
cosLookup[14234] <= 0.20459053;
cosLookup[14235] <= 0.204496678;
cosLookup[14236] <= 0.204402823;
cosLookup[14237] <= 0.204308967;
cosLookup[14238] <= 0.204215109;
cosLookup[14239] <= 0.204121249;
cosLookup[14240] <= 0.204027387;
cosLookup[14241] <= 0.203933523;
cosLookup[14242] <= 0.203839657;
cosLookup[14243] <= 0.20374579;
cosLookup[14244] <= 0.20365192;
cosLookup[14245] <= 0.203558049;
cosLookup[14246] <= 0.203464176;
cosLookup[14247] <= 0.203370301;
cosLookup[14248] <= 0.203276424;
cosLookup[14249] <= 0.203182545;
cosLookup[14250] <= 0.203088665;
cosLookup[14251] <= 0.202994782;
cosLookup[14252] <= 0.202900898;
cosLookup[14253] <= 0.202807012;
cosLookup[14254] <= 0.202713124;
cosLookup[14255] <= 0.202619234;
cosLookup[14256] <= 0.202525342;
cosLookup[14257] <= 0.202431448;
cosLookup[14258] <= 0.202337553;
cosLookup[14259] <= 0.202243655;
cosLookup[14260] <= 0.202149756;
cosLookup[14261] <= 0.202055855;
cosLookup[14262] <= 0.201961952;
cosLookup[14263] <= 0.201868047;
cosLookup[14264] <= 0.20177414;
cosLookup[14265] <= 0.201680232;
cosLookup[14266] <= 0.201586322;
cosLookup[14267] <= 0.201492409;
cosLookup[14268] <= 0.201398495;
cosLookup[14269] <= 0.201304579;
cosLookup[14270] <= 0.201210661;
cosLookup[14271] <= 0.201116742;
cosLookup[14272] <= 0.20102282;
cosLookup[14273] <= 0.200928897;
cosLookup[14274] <= 0.200834972;
cosLookup[14275] <= 0.200741045;
cosLookup[14276] <= 0.200647116;
cosLookup[14277] <= 0.200553185;
cosLookup[14278] <= 0.200459253;
cosLookup[14279] <= 0.200365318;
cosLookup[14280] <= 0.200271382;
cosLookup[14281] <= 0.200177444;
cosLookup[14282] <= 0.200083504;
cosLookup[14283] <= 0.199989562;
cosLookup[14284] <= 0.199895618;
cosLookup[14285] <= 0.199801673;
cosLookup[14286] <= 0.199707726;
cosLookup[14287] <= 0.199613777;
cosLookup[14288] <= 0.199519826;
cosLookup[14289] <= 0.199425873;
cosLookup[14290] <= 0.199331918;
cosLookup[14291] <= 0.199237962;
cosLookup[14292] <= 0.199144004;
cosLookup[14293] <= 0.199050043;
cosLookup[14294] <= 0.198956081;
cosLookup[14295] <= 0.198862118;
cosLookup[14296] <= 0.198768152;
cosLookup[14297] <= 0.198674185;
cosLookup[14298] <= 0.198580215;
cosLookup[14299] <= 0.198486244;
cosLookup[14300] <= 0.198392271;
cosLookup[14301] <= 0.198298297;
cosLookup[14302] <= 0.19820432;
cosLookup[14303] <= 0.198110342;
cosLookup[14304] <= 0.198016361;
cosLookup[14305] <= 0.197922379;
cosLookup[14306] <= 0.197828396;
cosLookup[14307] <= 0.19773441;
cosLookup[14308] <= 0.197640422;
cosLookup[14309] <= 0.197546433;
cosLookup[14310] <= 0.197452442;
cosLookup[14311] <= 0.197358449;
cosLookup[14312] <= 0.197264454;
cosLookup[14313] <= 0.197170458;
cosLookup[14314] <= 0.19707646;
cosLookup[14315] <= 0.196982459;
cosLookup[14316] <= 0.196888457;
cosLookup[14317] <= 0.196794454;
cosLookup[14318] <= 0.196700448;
cosLookup[14319] <= 0.196606441;
cosLookup[14320] <= 0.196512431;
cosLookup[14321] <= 0.19641842;
cosLookup[14322] <= 0.196324407;
cosLookup[14323] <= 0.196230393;
cosLookup[14324] <= 0.196136376;
cosLookup[14325] <= 0.196042358;
cosLookup[14326] <= 0.195948338;
cosLookup[14327] <= 0.195854316;
cosLookup[14328] <= 0.195760293;
cosLookup[14329] <= 0.195666267;
cosLookup[14330] <= 0.19557224;
cosLookup[14331] <= 0.195478211;
cosLookup[14332] <= 0.19538418;
cosLookup[14333] <= 0.195290147;
cosLookup[14334] <= 0.195196113;
cosLookup[14335] <= 0.195102077;
cosLookup[14336] <= 0.195008039;
cosLookup[14337] <= 0.194913999;
cosLookup[14338] <= 0.194819957;
cosLookup[14339] <= 0.194725914;
cosLookup[14340] <= 0.194631869;
cosLookup[14341] <= 0.194537822;
cosLookup[14342] <= 0.194443773;
cosLookup[14343] <= 0.194349722;
cosLookup[14344] <= 0.19425567;
cosLookup[14345] <= 0.194161616;
cosLookup[14346] <= 0.19406756;
cosLookup[14347] <= 0.193973502;
cosLookup[14348] <= 0.193879443;
cosLookup[14349] <= 0.193785382;
cosLookup[14350] <= 0.193691318;
cosLookup[14351] <= 0.193597254;
cosLookup[14352] <= 0.193503187;
cosLookup[14353] <= 0.193409119;
cosLookup[14354] <= 0.193315049;
cosLookup[14355] <= 0.193220977;
cosLookup[14356] <= 0.193126903;
cosLookup[14357] <= 0.193032827;
cosLookup[14358] <= 0.19293875;
cosLookup[14359] <= 0.192844671;
cosLookup[14360] <= 0.19275059;
cosLookup[14361] <= 0.192656508;
cosLookup[14362] <= 0.192562423;
cosLookup[14363] <= 0.192468337;
cosLookup[14364] <= 0.192374249;
cosLookup[14365] <= 0.19228016;
cosLookup[14366] <= 0.192186068;
cosLookup[14367] <= 0.192091975;
cosLookup[14368] <= 0.19199788;
cosLookup[14369] <= 0.191903783;
cosLookup[14370] <= 0.191809685;
cosLookup[14371] <= 0.191715585;
cosLookup[14372] <= 0.191621483;
cosLookup[14373] <= 0.191527379;
cosLookup[14374] <= 0.191433273;
cosLookup[14375] <= 0.191339166;
cosLookup[14376] <= 0.191245057;
cosLookup[14377] <= 0.191150946;
cosLookup[14378] <= 0.191056834;
cosLookup[14379] <= 0.190962719;
cosLookup[14380] <= 0.190868603;
cosLookup[14381] <= 0.190774485;
cosLookup[14382] <= 0.190680366;
cosLookup[14383] <= 0.190586244;
cosLookup[14384] <= 0.190492121;
cosLookup[14385] <= 0.190397996;
cosLookup[14386] <= 0.19030387;
cosLookup[14387] <= 0.190209741;
cosLookup[14388] <= 0.190115611;
cosLookup[14389] <= 0.19002148;
cosLookup[14390] <= 0.189927346;
cosLookup[14391] <= 0.189833211;
cosLookup[14392] <= 0.189739074;
cosLookup[14393] <= 0.189644935;
cosLookup[14394] <= 0.189550794;
cosLookup[14395] <= 0.189456652;
cosLookup[14396] <= 0.189362508;
cosLookup[14397] <= 0.189268362;
cosLookup[14398] <= 0.189174214;
cosLookup[14399] <= 0.189080065;
cosLookup[14400] <= 0.188985914;
cosLookup[14401] <= 0.188891761;
cosLookup[14402] <= 0.188797607;
cosLookup[14403] <= 0.188703451;
cosLookup[14404] <= 0.188609293;
cosLookup[14405] <= 0.188515133;
cosLookup[14406] <= 0.188420972;
cosLookup[14407] <= 0.188326808;
cosLookup[14408] <= 0.188232644;
cosLookup[14409] <= 0.188138477;
cosLookup[14410] <= 0.188044309;
cosLookup[14411] <= 0.187950139;
cosLookup[14412] <= 0.187855967;
cosLookup[14413] <= 0.187761793;
cosLookup[14414] <= 0.187667618;
cosLookup[14415] <= 0.187573441;
cosLookup[14416] <= 0.187479262;
cosLookup[14417] <= 0.187385082;
cosLookup[14418] <= 0.1872909;
cosLookup[14419] <= 0.187196716;
cosLookup[14420] <= 0.18710253;
cosLookup[14421] <= 0.187008343;
cosLookup[14422] <= 0.186914154;
cosLookup[14423] <= 0.186819963;
cosLookup[14424] <= 0.186725771;
cosLookup[14425] <= 0.186631576;
cosLookup[14426] <= 0.186537381;
cosLookup[14427] <= 0.186443183;
cosLookup[14428] <= 0.186348984;
cosLookup[14429] <= 0.186254783;
cosLookup[14430] <= 0.18616058;
cosLookup[14431] <= 0.186066375;
cosLookup[14432] <= 0.185972169;
cosLookup[14433] <= 0.185877961;
cosLookup[14434] <= 0.185783752;
cosLookup[14435] <= 0.18568954;
cosLookup[14436] <= 0.185595327;
cosLookup[14437] <= 0.185501113;
cosLookup[14438] <= 0.185406896;
cosLookup[14439] <= 0.185312678;
cosLookup[14440] <= 0.185218458;
cosLookup[14441] <= 0.185124237;
cosLookup[14442] <= 0.185030014;
cosLookup[14443] <= 0.184935789;
cosLookup[14444] <= 0.184841562;
cosLookup[14445] <= 0.184747334;
cosLookup[14446] <= 0.184653104;
cosLookup[14447] <= 0.184558872;
cosLookup[14448] <= 0.184464638;
cosLookup[14449] <= 0.184370403;
cosLookup[14450] <= 0.184276166;
cosLookup[14451] <= 0.184181928;
cosLookup[14452] <= 0.184087688;
cosLookup[14453] <= 0.183993446;
cosLookup[14454] <= 0.183899202;
cosLookup[14455] <= 0.183804957;
cosLookup[14456] <= 0.18371071;
cosLookup[14457] <= 0.183616461;
cosLookup[14458] <= 0.183522211;
cosLookup[14459] <= 0.183427959;
cosLookup[14460] <= 0.183333705;
cosLookup[14461] <= 0.18323945;
cosLookup[14462] <= 0.183145193;
cosLookup[14463] <= 0.183050934;
cosLookup[14464] <= 0.182956674;
cosLookup[14465] <= 0.182862411;
cosLookup[14466] <= 0.182768148;
cosLookup[14467] <= 0.182673882;
cosLookup[14468] <= 0.182579615;
cosLookup[14469] <= 0.182485346;
cosLookup[14470] <= 0.182391076;
cosLookup[14471] <= 0.182296803;
cosLookup[14472] <= 0.182202529;
cosLookup[14473] <= 0.182108254;
cosLookup[14474] <= 0.182013977;
cosLookup[14475] <= 0.181919698;
cosLookup[14476] <= 0.181825417;
cosLookup[14477] <= 0.181731135;
cosLookup[14478] <= 0.181636851;
cosLookup[14479] <= 0.181542565;
cosLookup[14480] <= 0.181448278;
cosLookup[14481] <= 0.181353989;
cosLookup[14482] <= 0.181259699;
cosLookup[14483] <= 0.181165406;
cosLookup[14484] <= 0.181071112;
cosLookup[14485] <= 0.180976817;
cosLookup[14486] <= 0.18088252;
cosLookup[14487] <= 0.180788221;
cosLookup[14488] <= 0.18069392;
cosLookup[14489] <= 0.180599618;
cosLookup[14490] <= 0.180505314;
cosLookup[14491] <= 0.180411008;
cosLookup[14492] <= 0.180316701;
cosLookup[14493] <= 0.180222392;
cosLookup[14494] <= 0.180128082;
cosLookup[14495] <= 0.18003377;
cosLookup[14496] <= 0.179939456;
cosLookup[14497] <= 0.17984514;
cosLookup[14498] <= 0.179750823;
cosLookup[14499] <= 0.179656504;
cosLookup[14500] <= 0.179562184;
cosLookup[14501] <= 0.179467862;
cosLookup[14502] <= 0.179373538;
cosLookup[14503] <= 0.179279212;
cosLookup[14504] <= 0.179184885;
cosLookup[14505] <= 0.179090557;
cosLookup[14506] <= 0.178996226;
cosLookup[14507] <= 0.178901894;
cosLookup[14508] <= 0.178807561;
cosLookup[14509] <= 0.178713225;
cosLookup[14510] <= 0.178618889;
cosLookup[14511] <= 0.17852455;
cosLookup[14512] <= 0.17843021;
cosLookup[14513] <= 0.178335868;
cosLookup[14514] <= 0.178241524;
cosLookup[14515] <= 0.178147179;
cosLookup[14516] <= 0.178052833;
cosLookup[14517] <= 0.177958484;
cosLookup[14518] <= 0.177864134;
cosLookup[14519] <= 0.177769782;
cosLookup[14520] <= 0.177675429;
cosLookup[14521] <= 0.177581074;
cosLookup[14522] <= 0.177486718;
cosLookup[14523] <= 0.177392359;
cosLookup[14524] <= 0.177298;
cosLookup[14525] <= 0.177203638;
cosLookup[14526] <= 0.177109275;
cosLookup[14527] <= 0.17701491;
cosLookup[14528] <= 0.176920544;
cosLookup[14529] <= 0.176826176;
cosLookup[14530] <= 0.176731806;
cosLookup[14531] <= 0.176637435;
cosLookup[14532] <= 0.176543062;
cosLookup[14533] <= 0.176448688;
cosLookup[14534] <= 0.176354312;
cosLookup[14535] <= 0.176259934;
cosLookup[14536] <= 0.176165555;
cosLookup[14537] <= 0.176071174;
cosLookup[14538] <= 0.175976791;
cosLookup[14539] <= 0.175882407;
cosLookup[14540] <= 0.175788021;
cosLookup[14541] <= 0.175693634;
cosLookup[14542] <= 0.175599245;
cosLookup[14543] <= 0.175504854;
cosLookup[14544] <= 0.175410462;
cosLookup[14545] <= 0.175316068;
cosLookup[14546] <= 0.175221672;
cosLookup[14547] <= 0.175127275;
cosLookup[14548] <= 0.175032877;
cosLookup[14549] <= 0.174938476;
cosLookup[14550] <= 0.174844074;
cosLookup[14551] <= 0.174749671;
cosLookup[14552] <= 0.174655266;
cosLookup[14553] <= 0.174560859;
cosLookup[14554] <= 0.17446645;
cosLookup[14555] <= 0.174372041;
cosLookup[14556] <= 0.174277629;
cosLookup[14557] <= 0.174183216;
cosLookup[14558] <= 0.174088801;
cosLookup[14559] <= 0.173994385;
cosLookup[14560] <= 0.173899967;
cosLookup[14561] <= 0.173805547;
cosLookup[14562] <= 0.173711126;
cosLookup[14563] <= 0.173616703;
cosLookup[14564] <= 0.173522279;
cosLookup[14565] <= 0.173427853;
cosLookup[14566] <= 0.173333425;
cosLookup[14567] <= 0.173238996;
cosLookup[14568] <= 0.173144566;
cosLookup[14569] <= 0.173050133;
cosLookup[14570] <= 0.172955699;
cosLookup[14571] <= 0.172861264;
cosLookup[14572] <= 0.172766827;
cosLookup[14573] <= 0.172672388;
cosLookup[14574] <= 0.172577948;
cosLookup[14575] <= 0.172483506;
cosLookup[14576] <= 0.172389062;
cosLookup[14577] <= 0.172294617;
cosLookup[14578] <= 0.172200171;
cosLookup[14579] <= 0.172105723;
cosLookup[14580] <= 0.172011273;
cosLookup[14581] <= 0.171916822;
cosLookup[14582] <= 0.171822369;
cosLookup[14583] <= 0.171727914;
cosLookup[14584] <= 0.171633458;
cosLookup[14585] <= 0.171539;
cosLookup[14586] <= 0.171444541;
cosLookup[14587] <= 0.17135008;
cosLookup[14588] <= 0.171255618;
cosLookup[14589] <= 0.171161154;
cosLookup[14590] <= 0.171066688;
cosLookup[14591] <= 0.170972221;
cosLookup[14592] <= 0.170877753;
cosLookup[14593] <= 0.170783282;
cosLookup[14594] <= 0.17068881;
cosLookup[14595] <= 0.170594337;
cosLookup[14596] <= 0.170499862;
cosLookup[14597] <= 0.170405386;
cosLookup[14598] <= 0.170310907;
cosLookup[14599] <= 0.170216428;
cosLookup[14600] <= 0.170121947;
cosLookup[14601] <= 0.170027464;
cosLookup[14602] <= 0.169932979;
cosLookup[14603] <= 0.169838493;
cosLookup[14604] <= 0.169744006;
cosLookup[14605] <= 0.169649517;
cosLookup[14606] <= 0.169555026;
cosLookup[14607] <= 0.169460534;
cosLookup[14608] <= 0.16936604;
cosLookup[14609] <= 0.169271545;
cosLookup[14610] <= 0.169177048;
cosLookup[14611] <= 0.16908255;
cosLookup[14612] <= 0.16898805;
cosLookup[14613] <= 0.168893548;
cosLookup[14614] <= 0.168799045;
cosLookup[14615] <= 0.168704541;
cosLookup[14616] <= 0.168610035;
cosLookup[14617] <= 0.168515527;
cosLookup[14618] <= 0.168421018;
cosLookup[14619] <= 0.168326507;
cosLookup[14620] <= 0.168231995;
cosLookup[14621] <= 0.168137481;
cosLookup[14622] <= 0.168042965;
cosLookup[14623] <= 0.167948448;
cosLookup[14624] <= 0.16785393;
cosLookup[14625] <= 0.16775941;
cosLookup[14626] <= 0.167664888;
cosLookup[14627] <= 0.167570365;
cosLookup[14628] <= 0.16747584;
cosLookup[14629] <= 0.167381314;
cosLookup[14630] <= 0.167286786;
cosLookup[14631] <= 0.167192257;
cosLookup[14632] <= 0.167097726;
cosLookup[14633] <= 0.167003194;
cosLookup[14634] <= 0.16690866;
cosLookup[14635] <= 0.166814124;
cosLookup[14636] <= 0.166719587;
cosLookup[14637] <= 0.166625049;
cosLookup[14638] <= 0.166530509;
cosLookup[14639] <= 0.166435967;
cosLookup[14640] <= 0.166341424;
cosLookup[14641] <= 0.166246879;
cosLookup[14642] <= 0.166152333;
cosLookup[14643] <= 0.166057786;
cosLookup[14644] <= 0.165963236;
cosLookup[14645] <= 0.165868686;
cosLookup[14646] <= 0.165774133;
cosLookup[14647] <= 0.165679579;
cosLookup[14648] <= 0.165585024;
cosLookup[14649] <= 0.165490467;
cosLookup[14650] <= 0.165395909;
cosLookup[14651] <= 0.165301349;
cosLookup[14652] <= 0.165206788;
cosLookup[14653] <= 0.165112225;
cosLookup[14654] <= 0.16501766;
cosLookup[14655] <= 0.164923094;
cosLookup[14656] <= 0.164828527;
cosLookup[14657] <= 0.164733958;
cosLookup[14658] <= 0.164639387;
cosLookup[14659] <= 0.164544815;
cosLookup[14660] <= 0.164450242;
cosLookup[14661] <= 0.164355667;
cosLookup[14662] <= 0.16426109;
cosLookup[14663] <= 0.164166512;
cosLookup[14664] <= 0.164071933;
cosLookup[14665] <= 0.163977352;
cosLookup[14666] <= 0.163882769;
cosLookup[14667] <= 0.163788185;
cosLookup[14668] <= 0.163693599;
cosLookup[14669] <= 0.163599012;
cosLookup[14670] <= 0.163504424;
cosLookup[14671] <= 0.163409833;
cosLookup[14672] <= 0.163315242;
cosLookup[14673] <= 0.163220649;
cosLookup[14674] <= 0.163126054;
cosLookup[14675] <= 0.163031458;
cosLookup[14676] <= 0.16293686;
cosLookup[14677] <= 0.162842261;
cosLookup[14678] <= 0.162747661;
cosLookup[14679] <= 0.162653058;
cosLookup[14680] <= 0.162558455;
cosLookup[14681] <= 0.16246385;
cosLookup[14682] <= 0.162369243;
cosLookup[14683] <= 0.162274635;
cosLookup[14684] <= 0.162180026;
cosLookup[14685] <= 0.162085414;
cosLookup[14686] <= 0.161990802;
cosLookup[14687] <= 0.161896188;
cosLookup[14688] <= 0.161801572;
cosLookup[14689] <= 0.161706955;
cosLookup[14690] <= 0.161612337;
cosLookup[14691] <= 0.161517717;
cosLookup[14692] <= 0.161423095;
cosLookup[14693] <= 0.161328472;
cosLookup[14694] <= 0.161233848;
cosLookup[14695] <= 0.161139222;
cosLookup[14696] <= 0.161044595;
cosLookup[14697] <= 0.160949966;
cosLookup[14698] <= 0.160855335;
cosLookup[14699] <= 0.160760704;
cosLookup[14700] <= 0.16066607;
cosLookup[14701] <= 0.160571435;
cosLookup[14702] <= 0.160476799;
cosLookup[14703] <= 0.160382161;
cosLookup[14704] <= 0.160287522;
cosLookup[14705] <= 0.160192881;
cosLookup[14706] <= 0.160098239;
cosLookup[14707] <= 0.160003596;
cosLookup[14708] <= 0.159908951;
cosLookup[14709] <= 0.159814304;
cosLookup[14710] <= 0.159719656;
cosLookup[14711] <= 0.159625006;
cosLookup[14712] <= 0.159530355;
cosLookup[14713] <= 0.159435703;
cosLookup[14714] <= 0.159341049;
cosLookup[14715] <= 0.159246394;
cosLookup[14716] <= 0.159151737;
cosLookup[14717] <= 0.159057078;
cosLookup[14718] <= 0.158962419;
cosLookup[14719] <= 0.158867757;
cosLookup[14720] <= 0.158773095;
cosLookup[14721] <= 0.158678431;
cosLookup[14722] <= 0.158583765;
cosLookup[14723] <= 0.158489098;
cosLookup[14724] <= 0.158394429;
cosLookup[14725] <= 0.158299759;
cosLookup[14726] <= 0.158205088;
cosLookup[14727] <= 0.158110415;
cosLookup[14728] <= 0.158015741;
cosLookup[14729] <= 0.157921065;
cosLookup[14730] <= 0.157826388;
cosLookup[14731] <= 0.157731709;
cosLookup[14732] <= 0.157637029;
cosLookup[14733] <= 0.157542347;
cosLookup[14734] <= 0.157447664;
cosLookup[14735] <= 0.15735298;
cosLookup[14736] <= 0.157258294;
cosLookup[14737] <= 0.157163606;
cosLookup[14738] <= 0.157068917;
cosLookup[14739] <= 0.156974227;
cosLookup[14740] <= 0.156879535;
cosLookup[14741] <= 0.156784842;
cosLookup[14742] <= 0.156690148;
cosLookup[14743] <= 0.156595452;
cosLookup[14744] <= 0.156500754;
cosLookup[14745] <= 0.156406055;
cosLookup[14746] <= 0.156311355;
cosLookup[14747] <= 0.156216653;
cosLookup[14748] <= 0.15612195;
cosLookup[14749] <= 0.156027245;
cosLookup[14750] <= 0.155932539;
cosLookup[14751] <= 0.155837831;
cosLookup[14752] <= 0.155743123;
cosLookup[14753] <= 0.155648412;
cosLookup[14754] <= 0.1555537;
cosLookup[14755] <= 0.155458987;
cosLookup[14756] <= 0.155364272;
cosLookup[14757] <= 0.155269556;
cosLookup[14758] <= 0.155174839;
cosLookup[14759] <= 0.15508012;
cosLookup[14760] <= 0.154985399;
cosLookup[14761] <= 0.154890677;
cosLookup[14762] <= 0.154795954;
cosLookup[14763] <= 0.15470123;
cosLookup[14764] <= 0.154606503;
cosLookup[14765] <= 0.154511776;
cosLookup[14766] <= 0.154417047;
cosLookup[14767] <= 0.154322317;
cosLookup[14768] <= 0.154227585;
cosLookup[14769] <= 0.154132852;
cosLookup[14770] <= 0.154038117;
cosLookup[14771] <= 0.153943381;
cosLookup[14772] <= 0.153848644;
cosLookup[14773] <= 0.153753905;
cosLookup[14774] <= 0.153659164;
cosLookup[14775] <= 0.153564423;
cosLookup[14776] <= 0.15346968;
cosLookup[14777] <= 0.153374935;
cosLookup[14778] <= 0.153280189;
cosLookup[14779] <= 0.153185442;
cosLookup[14780] <= 0.153090693;
cosLookup[14781] <= 0.152995943;
cosLookup[14782] <= 0.152901192;
cosLookup[14783] <= 0.152806439;
cosLookup[14784] <= 0.152711684;
cosLookup[14785] <= 0.152616928;
cosLookup[14786] <= 0.152522171;
cosLookup[14787] <= 0.152427413;
cosLookup[14788] <= 0.152332653;
cosLookup[14789] <= 0.152237891;
cosLookup[14790] <= 0.152143129;
cosLookup[14791] <= 0.152048364;
cosLookup[14792] <= 0.151953599;
cosLookup[14793] <= 0.151858832;
cosLookup[14794] <= 0.151764064;
cosLookup[14795] <= 0.151669294;
cosLookup[14796] <= 0.151574523;
cosLookup[14797] <= 0.15147975;
cosLookup[14798] <= 0.151384976;
cosLookup[14799] <= 0.151290201;
cosLookup[14800] <= 0.151195424;
cosLookup[14801] <= 0.151100646;
cosLookup[14802] <= 0.151005867;
cosLookup[14803] <= 0.150911086;
cosLookup[14804] <= 0.150816303;
cosLookup[14805] <= 0.15072152;
cosLookup[14806] <= 0.150626735;
cosLookup[14807] <= 0.150531948;
cosLookup[14808] <= 0.15043716;
cosLookup[14809] <= 0.150342371;
cosLookup[14810] <= 0.150247581;
cosLookup[14811] <= 0.150152789;
cosLookup[14812] <= 0.150057995;
cosLookup[14813] <= 0.149963201;
cosLookup[14814] <= 0.149868405;
cosLookup[14815] <= 0.149773607;
cosLookup[14816] <= 0.149678808;
cosLookup[14817] <= 0.149584008;
cosLookup[14818] <= 0.149489206;
cosLookup[14819] <= 0.149394404;
cosLookup[14820] <= 0.149299599;
cosLookup[14821] <= 0.149204793;
cosLookup[14822] <= 0.149109986;
cosLookup[14823] <= 0.149015178;
cosLookup[14824] <= 0.148920368;
cosLookup[14825] <= 0.148825557;
cosLookup[14826] <= 0.148730744;
cosLookup[14827] <= 0.14863593;
cosLookup[14828] <= 0.148541115;
cosLookup[14829] <= 0.148446298;
cosLookup[14830] <= 0.14835148;
cosLookup[14831] <= 0.148256661;
cosLookup[14832] <= 0.14816184;
cosLookup[14833] <= 0.148067018;
cosLookup[14834] <= 0.147972195;
cosLookup[14835] <= 0.14787737;
cosLookup[14836] <= 0.147782544;
cosLookup[14837] <= 0.147687716;
cosLookup[14838] <= 0.147592887;
cosLookup[14839] <= 0.147498057;
cosLookup[14840] <= 0.147403225;
cosLookup[14841] <= 0.147308392;
cosLookup[14842] <= 0.147213558;
cosLookup[14843] <= 0.147118722;
cosLookup[14844] <= 0.147023885;
cosLookup[14845] <= 0.146929047;
cosLookup[14846] <= 0.146834207;
cosLookup[14847] <= 0.146739366;
cosLookup[14848] <= 0.146644523;
cosLookup[14849] <= 0.14654968;
cosLookup[14850] <= 0.146454834;
cosLookup[14851] <= 0.146359988;
cosLookup[14852] <= 0.14626514;
cosLookup[14853] <= 0.146170291;
cosLookup[14854] <= 0.14607544;
cosLookup[14855] <= 0.145980589;
cosLookup[14856] <= 0.145885735;
cosLookup[14857] <= 0.145790881;
cosLookup[14858] <= 0.145696025;
cosLookup[14859] <= 0.145601168;
cosLookup[14860] <= 0.145506309;
cosLookup[14861] <= 0.145411449;
cosLookup[14862] <= 0.145316588;
cosLookup[14863] <= 0.145221725;
cosLookup[14864] <= 0.145126862;
cosLookup[14865] <= 0.145031996;
cosLookup[14866] <= 0.14493713;
cosLookup[14867] <= 0.144842262;
cosLookup[14868] <= 0.144747393;
cosLookup[14869] <= 0.144652522;
cosLookup[14870] <= 0.14455765;
cosLookup[14871] <= 0.144462777;
cosLookup[14872] <= 0.144367902;
cosLookup[14873] <= 0.144273026;
cosLookup[14874] <= 0.144178149;
cosLookup[14875] <= 0.144083271;
cosLookup[14876] <= 0.143988391;
cosLookup[14877] <= 0.14389351;
cosLookup[14878] <= 0.143798627;
cosLookup[14879] <= 0.143703743;
cosLookup[14880] <= 0.143608858;
cosLookup[14881] <= 0.143513972;
cosLookup[14882] <= 0.143419084;
cosLookup[14883] <= 0.143324195;
cosLookup[14884] <= 0.143229304;
cosLookup[14885] <= 0.143134413;
cosLookup[14886] <= 0.143039519;
cosLookup[14887] <= 0.142944625;
cosLookup[14888] <= 0.142849729;
cosLookup[14889] <= 0.142754832;
cosLookup[14890] <= 0.142659934;
cosLookup[14891] <= 0.142565034;
cosLookup[14892] <= 0.142470134;
cosLookup[14893] <= 0.142375231;
cosLookup[14894] <= 0.142280328;
cosLookup[14895] <= 0.142185423;
cosLookup[14896] <= 0.142090517;
cosLookup[14897] <= 0.141995609;
cosLookup[14898] <= 0.1419007;
cosLookup[14899] <= 0.14180579;
cosLookup[14900] <= 0.141710879;
cosLookup[14901] <= 0.141615966;
cosLookup[14902] <= 0.141521052;
cosLookup[14903] <= 0.141426137;
cosLookup[14904] <= 0.14133122;
cosLookup[14905] <= 0.141236302;
cosLookup[14906] <= 0.141141383;
cosLookup[14907] <= 0.141046463;
cosLookup[14908] <= 0.140951541;
cosLookup[14909] <= 0.140856618;
cosLookup[14910] <= 0.140761694;
cosLookup[14911] <= 0.140666768;
cosLookup[14912] <= 0.140571841;
cosLookup[14913] <= 0.140476913;
cosLookup[14914] <= 0.140381983;
cosLookup[14915] <= 0.140287052;
cosLookup[14916] <= 0.14019212;
cosLookup[14917] <= 0.140097187;
cosLookup[14918] <= 0.140002252;
cosLookup[14919] <= 0.139907316;
cosLookup[14920] <= 0.139812379;
cosLookup[14921] <= 0.13971744;
cosLookup[14922] <= 0.1396225;
cosLookup[14923] <= 0.139527559;
cosLookup[14924] <= 0.139432617;
cosLookup[14925] <= 0.139337673;
cosLookup[14926] <= 0.139242728;
cosLookup[14927] <= 0.139147782;
cosLookup[14928] <= 0.139052834;
cosLookup[14929] <= 0.138957885;
cosLookup[14930] <= 0.138862935;
cosLookup[14931] <= 0.138767984;
cosLookup[14932] <= 0.138673031;
cosLookup[14933] <= 0.138578077;
cosLookup[14934] <= 0.138483122;
cosLookup[14935] <= 0.138388166;
cosLookup[14936] <= 0.138293208;
cosLookup[14937] <= 0.138198249;
cosLookup[14938] <= 0.138103289;
cosLookup[14939] <= 0.138008327;
cosLookup[14940] <= 0.137913364;
cosLookup[14941] <= 0.1378184;
cosLookup[14942] <= 0.137723435;
cosLookup[14943] <= 0.137628468;
cosLookup[14944] <= 0.1375335;
cosLookup[14945] <= 0.137438531;
cosLookup[14946] <= 0.137343561;
cosLookup[14947] <= 0.137248589;
cosLookup[14948] <= 0.137153616;
cosLookup[14949] <= 0.137058642;
cosLookup[14950] <= 0.136963667;
cosLookup[14951] <= 0.13686869;
cosLookup[14952] <= 0.136773712;
cosLookup[14953] <= 0.136678733;
cosLookup[14954] <= 0.136583752;
cosLookup[14955] <= 0.13648877;
cosLookup[14956] <= 0.136393787;
cosLookup[14957] <= 0.136298803;
cosLookup[14958] <= 0.136203818;
cosLookup[14959] <= 0.136108831;
cosLookup[14960] <= 0.136013843;
cosLookup[14961] <= 0.135918854;
cosLookup[14962] <= 0.135823863;
cosLookup[14963] <= 0.135728871;
cosLookup[14964] <= 0.135633878;
cosLookup[14965] <= 0.135538884;
cosLookup[14966] <= 0.135443889;
cosLookup[14967] <= 0.135348892;
cosLookup[14968] <= 0.135253894;
cosLookup[14969] <= 0.135158895;
cosLookup[14970] <= 0.135063894;
cosLookup[14971] <= 0.134968892;
cosLookup[14972] <= 0.13487389;
cosLookup[14973] <= 0.134778885;
cosLookup[14974] <= 0.13468388;
cosLookup[14975] <= 0.134588873;
cosLookup[14976] <= 0.134493865;
cosLookup[14977] <= 0.134398856;
cosLookup[14978] <= 0.134303846;
cosLookup[14979] <= 0.134208834;
cosLookup[14980] <= 0.134113821;
cosLookup[14981] <= 0.134018807;
cosLookup[14982] <= 0.133923792;
cosLookup[14983] <= 0.133828775;
cosLookup[14984] <= 0.133733758;
cosLookup[14985] <= 0.133638739;
cosLookup[14986] <= 0.133543718;
cosLookup[14987] <= 0.133448697;
cosLookup[14988] <= 0.133353674;
cosLookup[14989] <= 0.13325865;
cosLookup[14990] <= 0.133163625;
cosLookup[14991] <= 0.133068599;
cosLookup[14992] <= 0.132973571;
cosLookup[14993] <= 0.132878542;
cosLookup[14994] <= 0.132783512;
cosLookup[14995] <= 0.132688481;
cosLookup[14996] <= 0.132593449;
cosLookup[14997] <= 0.132498415;
cosLookup[14998] <= 0.13240338;
cosLookup[14999] <= 0.132308344;
cosLookup[15000] <= 0.132213307;
cosLookup[15001] <= 0.132118268;
cosLookup[15002] <= 0.132023228;
cosLookup[15003] <= 0.131928187;
cosLookup[15004] <= 0.131833145;
cosLookup[15005] <= 0.131738102;
cosLookup[15006] <= 0.131643057;
cosLookup[15007] <= 0.131548011;
cosLookup[15008] <= 0.131452964;
cosLookup[15009] <= 0.131357916;
cosLookup[15010] <= 0.131262866;
cosLookup[15011] <= 0.131167816;
cosLookup[15012] <= 0.131072764;
cosLookup[15013] <= 0.130977711;
cosLookup[15014] <= 0.130882656;
cosLookup[15015] <= 0.130787601;
cosLookup[15016] <= 0.130692544;
cosLookup[15017] <= 0.130597486;
cosLookup[15018] <= 0.130502427;
cosLookup[15019] <= 0.130407367;
cosLookup[15020] <= 0.130312306;
cosLookup[15021] <= 0.130217243;
cosLookup[15022] <= 0.130122179;
cosLookup[15023] <= 0.130027114;
cosLookup[15024] <= 0.129932048;
cosLookup[15025] <= 0.12983698;
cosLookup[15026] <= 0.129741912;
cosLookup[15027] <= 0.129646842;
cosLookup[15028] <= 0.129551771;
cosLookup[15029] <= 0.129456698;
cosLookup[15030] <= 0.129361625;
cosLookup[15031] <= 0.12926655;
cosLookup[15032] <= 0.129171475;
cosLookup[15033] <= 0.129076398;
cosLookup[15034] <= 0.128981319;
cosLookup[15035] <= 0.12888624;
cosLookup[15036] <= 0.128791159;
cosLookup[15037] <= 0.128696078;
cosLookup[15038] <= 0.128600995;
cosLookup[15039] <= 0.128505911;
cosLookup[15040] <= 0.128410825;
cosLookup[15041] <= 0.128315739;
cosLookup[15042] <= 0.128220651;
cosLookup[15043] <= 0.128125563;
cosLookup[15044] <= 0.128030473;
cosLookup[15045] <= 0.127935381;
cosLookup[15046] <= 0.127840289;
cosLookup[15047] <= 0.127745195;
cosLookup[15048] <= 0.127650101;
cosLookup[15049] <= 0.127555005;
cosLookup[15050] <= 0.127459908;
cosLookup[15051] <= 0.12736481;
cosLookup[15052] <= 0.12726971;
cosLookup[15053] <= 0.12717461;
cosLookup[15054] <= 0.127079508;
cosLookup[15055] <= 0.126984405;
cosLookup[15056] <= 0.126889301;
cosLookup[15057] <= 0.126794196;
cosLookup[15058] <= 0.126699089;
cosLookup[15059] <= 0.126603982;
cosLookup[15060] <= 0.126508873;
cosLookup[15061] <= 0.126413763;
cosLookup[15062] <= 0.126318652;
cosLookup[15063] <= 0.12622354;
cosLookup[15064] <= 0.126128427;
cosLookup[15065] <= 0.126033312;
cosLookup[15066] <= 0.125938196;
cosLookup[15067] <= 0.12584308;
cosLookup[15068] <= 0.125747962;
cosLookup[15069] <= 0.125652842;
cosLookup[15070] <= 0.125557722;
cosLookup[15071] <= 0.125462601;
cosLookup[15072] <= 0.125367478;
cosLookup[15073] <= 0.125272354;
cosLookup[15074] <= 0.125177229;
cosLookup[15075] <= 0.125082103;
cosLookup[15076] <= 0.124986976;
cosLookup[15077] <= 0.124891848;
cosLookup[15078] <= 0.124796718;
cosLookup[15079] <= 0.124701587;
cosLookup[15080] <= 0.124606456;
cosLookup[15081] <= 0.124511323;
cosLookup[15082] <= 0.124416189;
cosLookup[15083] <= 0.124321053;
cosLookup[15084] <= 0.124225917;
cosLookup[15085] <= 0.124130779;
cosLookup[15086] <= 0.124035641;
cosLookup[15087] <= 0.123940501;
cosLookup[15088] <= 0.12384536;
cosLookup[15089] <= 0.123750218;
cosLookup[15090] <= 0.123655075;
cosLookup[15091] <= 0.12355993;
cosLookup[15092] <= 0.123464785;
cosLookup[15093] <= 0.123369638;
cosLookup[15094] <= 0.12327449;
cosLookup[15095] <= 0.123179341;
cosLookup[15096] <= 0.123084191;
cosLookup[15097] <= 0.12298904;
cosLookup[15098] <= 0.122893888;
cosLookup[15099] <= 0.122798734;
cosLookup[15100] <= 0.12270358;
cosLookup[15101] <= 0.122608424;
cosLookup[15102] <= 0.122513267;
cosLookup[15103] <= 0.122418109;
cosLookup[15104] <= 0.12232295;
cosLookup[15105] <= 0.12222779;
cosLookup[15106] <= 0.122132629;
cosLookup[15107] <= 0.122037466;
cosLookup[15108] <= 0.121942303;
cosLookup[15109] <= 0.121847138;
cosLookup[15110] <= 0.121751972;
cosLookup[15111] <= 0.121656805;
cosLookup[15112] <= 0.121561637;
cosLookup[15113] <= 0.121466468;
cosLookup[15114] <= 0.121371298;
cosLookup[15115] <= 0.121276127;
cosLookup[15116] <= 0.121180954;
cosLookup[15117] <= 0.121085781;
cosLookup[15118] <= 0.120990606;
cosLookup[15119] <= 0.12089543;
cosLookup[15120] <= 0.120800253;
cosLookup[15121] <= 0.120705075;
cosLookup[15122] <= 0.120609896;
cosLookup[15123] <= 0.120514715;
cosLookup[15124] <= 0.120419534;
cosLookup[15125] <= 0.120324352;
cosLookup[15126] <= 0.120229168;
cosLookup[15127] <= 0.120133983;
cosLookup[15128] <= 0.120038797;
cosLookup[15129] <= 0.119943611;
cosLookup[15130] <= 0.119848423;
cosLookup[15131] <= 0.119753233;
cosLookup[15132] <= 0.119658043;
cosLookup[15133] <= 0.119562852;
cosLookup[15134] <= 0.119467659;
cosLookup[15135] <= 0.119372466;
cosLookup[15136] <= 0.119277271;
cosLookup[15137] <= 0.119182076;
cosLookup[15138] <= 0.119086879;
cosLookup[15139] <= 0.118991681;
cosLookup[15140] <= 0.118896482;
cosLookup[15141] <= 0.118801282;
cosLookup[15142] <= 0.118706081;
cosLookup[15143] <= 0.118610878;
cosLookup[15144] <= 0.118515675;
cosLookup[15145] <= 0.118420471;
cosLookup[15146] <= 0.118325265;
cosLookup[15147] <= 0.118230058;
cosLookup[15148] <= 0.118134851;
cosLookup[15149] <= 0.118039642;
cosLookup[15150] <= 0.117944432;
cosLookup[15151] <= 0.117849221;
cosLookup[15152] <= 0.117754009;
cosLookup[15153] <= 0.117658796;
cosLookup[15154] <= 0.117563582;
cosLookup[15155] <= 0.117468366;
cosLookup[15156] <= 0.11737315;
cosLookup[15157] <= 0.117277932;
cosLookup[15158] <= 0.117182714;
cosLookup[15159] <= 0.117087494;
cosLookup[15160] <= 0.116992274;
cosLookup[15161] <= 0.116897052;
cosLookup[15162] <= 0.116801829;
cosLookup[15163] <= 0.116706605;
cosLookup[15164] <= 0.11661138;
cosLookup[15165] <= 0.116516154;
cosLookup[15166] <= 0.116420927;
cosLookup[15167] <= 0.116325699;
cosLookup[15168] <= 0.116230469;
cosLookup[15169] <= 0.116135239;
cosLookup[15170] <= 0.116040008;
cosLookup[15171] <= 0.115944775;
cosLookup[15172] <= 0.115849542;
cosLookup[15173] <= 0.115754307;
cosLookup[15174] <= 0.115659071;
cosLookup[15175] <= 0.115563835;
cosLookup[15176] <= 0.115468597;
cosLookup[15177] <= 0.115373358;
cosLookup[15178] <= 0.115278118;
cosLookup[15179] <= 0.115182877;
cosLookup[15180] <= 0.115087635;
cosLookup[15181] <= 0.114992392;
cosLookup[15182] <= 0.114897148;
cosLookup[15183] <= 0.114801903;
cosLookup[15184] <= 0.114706656;
cosLookup[15185] <= 0.114611409;
cosLookup[15186] <= 0.114516161;
cosLookup[15187] <= 0.114420911;
cosLookup[15188] <= 0.114325661;
cosLookup[15189] <= 0.114230409;
cosLookup[15190] <= 0.114135157;
cosLookup[15191] <= 0.114039903;
cosLookup[15192] <= 0.113944648;
cosLookup[15193] <= 0.113849393;
cosLookup[15194] <= 0.113754136;
cosLookup[15195] <= 0.113658878;
cosLookup[15196] <= 0.113563619;
cosLookup[15197] <= 0.113468359;
cosLookup[15198] <= 0.113373098;
cosLookup[15199] <= 0.113277836;
cosLookup[15200] <= 0.113182573;
cosLookup[15201] <= 0.113087309;
cosLookup[15202] <= 0.112992044;
cosLookup[15203] <= 0.112896778;
cosLookup[15204] <= 0.112801511;
cosLookup[15205] <= 0.112706243;
cosLookup[15206] <= 0.112610973;
cosLookup[15207] <= 0.112515703;
cosLookup[15208] <= 0.112420432;
cosLookup[15209] <= 0.112325159;
cosLookup[15210] <= 0.112229886;
cosLookup[15211] <= 0.112134612;
cosLookup[15212] <= 0.112039336;
cosLookup[15213] <= 0.11194406;
cosLookup[15214] <= 0.111848782;
cosLookup[15215] <= 0.111753504;
cosLookup[15216] <= 0.111658224;
cosLookup[15217] <= 0.111562943;
cosLookup[15218] <= 0.111467662;
cosLookup[15219] <= 0.111372379;
cosLookup[15220] <= 0.111277095;
cosLookup[15221] <= 0.111181811;
cosLookup[15222] <= 0.111086525;
cosLookup[15223] <= 0.110991238;
cosLookup[15224] <= 0.110895951;
cosLookup[15225] <= 0.110800662;
cosLookup[15226] <= 0.110705372;
cosLookup[15227] <= 0.110610081;
cosLookup[15228] <= 0.110514789;
cosLookup[15229] <= 0.110419496;
cosLookup[15230] <= 0.110324203;
cosLookup[15231] <= 0.110228908;
cosLookup[15232] <= 0.110133612;
cosLookup[15233] <= 0.110038315;
cosLookup[15234] <= 0.109943017;
cosLookup[15235] <= 0.109847718;
cosLookup[15236] <= 0.109752418;
cosLookup[15237] <= 0.109657117;
cosLookup[15238] <= 0.109561815;
cosLookup[15239] <= 0.109466512;
cosLookup[15240] <= 0.109371208;
cosLookup[15241] <= 0.109275903;
cosLookup[15242] <= 0.109180597;
cosLookup[15243] <= 0.10908529;
cosLookup[15244] <= 0.108989982;
cosLookup[15245] <= 0.108894673;
cosLookup[15246] <= 0.108799364;
cosLookup[15247] <= 0.108704053;
cosLookup[15248] <= 0.108608741;
cosLookup[15249] <= 0.108513428;
cosLookup[15250] <= 0.108418114;
cosLookup[15251] <= 0.108322799;
cosLookup[15252] <= 0.108227483;
cosLookup[15253] <= 0.108132166;
cosLookup[15254] <= 0.108036848;
cosLookup[15255] <= 0.107941529;
cosLookup[15256] <= 0.107846209;
cosLookup[15257] <= 0.107750888;
cosLookup[15258] <= 0.107655566;
cosLookup[15259] <= 0.107560243;
cosLookup[15260] <= 0.107464919;
cosLookup[15261] <= 0.107369594;
cosLookup[15262] <= 0.107274268;
cosLookup[15263] <= 0.107178941;
cosLookup[15264] <= 0.107083614;
cosLookup[15265] <= 0.106988285;
cosLookup[15266] <= 0.106892955;
cosLookup[15267] <= 0.106797624;
cosLookup[15268] <= 0.106702292;
cosLookup[15269] <= 0.10660696;
cosLookup[15270] <= 0.106511626;
cosLookup[15271] <= 0.106416291;
cosLookup[15272] <= 0.106320955;
cosLookup[15273] <= 0.106225619;
cosLookup[15274] <= 0.106130281;
cosLookup[15275] <= 0.106034942;
cosLookup[15276] <= 0.105939603;
cosLookup[15277] <= 0.105844262;
cosLookup[15278] <= 0.105748921;
cosLookup[15279] <= 0.105653578;
cosLookup[15280] <= 0.105558235;
cosLookup[15281] <= 0.10546289;
cosLookup[15282] <= 0.105367545;
cosLookup[15283] <= 0.105272198;
cosLookup[15284] <= 0.105176851;
cosLookup[15285] <= 0.105081503;
cosLookup[15286] <= 0.104986153;
cosLookup[15287] <= 0.104890803;
cosLookup[15288] <= 0.104795452;
cosLookup[15289] <= 0.1047001;
cosLookup[15290] <= 0.104604746;
cosLookup[15291] <= 0.104509392;
cosLookup[15292] <= 0.104414037;
cosLookup[15293] <= 0.104318681;
cosLookup[15294] <= 0.104223324;
cosLookup[15295] <= 0.104127966;
cosLookup[15296] <= 0.104032607;
cosLookup[15297] <= 0.103937247;
cosLookup[15298] <= 0.103841887;
cosLookup[15299] <= 0.103746525;
cosLookup[15300] <= 0.103651162;
cosLookup[15301] <= 0.103555798;
cosLookup[15302] <= 0.103460434;
cosLookup[15303] <= 0.103365068;
cosLookup[15304] <= 0.103269702;
cosLookup[15305] <= 0.103174334;
cosLookup[15306] <= 0.103078966;
cosLookup[15307] <= 0.102983596;
cosLookup[15308] <= 0.102888226;
cosLookup[15309] <= 0.102792855;
cosLookup[15310] <= 0.102697482;
cosLookup[15311] <= 0.102602109;
cosLookup[15312] <= 0.102506735;
cosLookup[15313] <= 0.10241136;
cosLookup[15314] <= 0.102315984;
cosLookup[15315] <= 0.102220607;
cosLookup[15316] <= 0.102125229;
cosLookup[15317] <= 0.10202985;
cosLookup[15318] <= 0.101934471;
cosLookup[15319] <= 0.10183909;
cosLookup[15320] <= 0.101743708;
cosLookup[15321] <= 0.101648326;
cosLookup[15322] <= 0.101552942;
cosLookup[15323] <= 0.101457558;
cosLookup[15324] <= 0.101362173;
cosLookup[15325] <= 0.101266786;
cosLookup[15326] <= 0.101171399;
cosLookup[15327] <= 0.101076011;
cosLookup[15328] <= 0.100980622;
cosLookup[15329] <= 0.100885232;
cosLookup[15330] <= 0.100789841;
cosLookup[15331] <= 0.100694449;
cosLookup[15332] <= 0.100599056;
cosLookup[15333] <= 0.100503662;
cosLookup[15334] <= 0.100408268;
cosLookup[15335] <= 0.100312872;
cosLookup[15336] <= 0.100217476;
cosLookup[15337] <= 0.100122078;
cosLookup[15338] <= 0.10002668;
cosLookup[15339] <= 0.099931281;
cosLookup[15340] <= 0.099835881;
cosLookup[15341] <= 0.099740479;
cosLookup[15342] <= 0.099645077;
cosLookup[15343] <= 0.099549675;
cosLookup[15344] <= 0.099454271;
cosLookup[15345] <= 0.099358866;
cosLookup[15346] <= 0.09926346;
cosLookup[15347] <= 0.099168054;
cosLookup[15348] <= 0.099072646;
cosLookup[15349] <= 0.098977238;
cosLookup[15350] <= 0.098881829;
cosLookup[15351] <= 0.098786418;
cosLookup[15352] <= 0.098691007;
cosLookup[15353] <= 0.098595595;
cosLookup[15354] <= 0.098500182;
cosLookup[15355] <= 0.098404768;
cosLookup[15356] <= 0.098309354;
cosLookup[15357] <= 0.098213938;
cosLookup[15358] <= 0.098118521;
cosLookup[15359] <= 0.098023104;
cosLookup[15360] <= 0.097927686;
cosLookup[15361] <= 0.097832266;
cosLookup[15362] <= 0.097736846;
cosLookup[15363] <= 0.097641425;
cosLookup[15364] <= 0.097546003;
cosLookup[15365] <= 0.09745058;
cosLookup[15366] <= 0.097355157;
cosLookup[15367] <= 0.097259732;
cosLookup[15368] <= 0.097164306;
cosLookup[15369] <= 0.09706888;
cosLookup[15370] <= 0.096973453;
cosLookup[15371] <= 0.096878024;
cosLookup[15372] <= 0.096782595;
cosLookup[15373] <= 0.096687165;
cosLookup[15374] <= 0.096591734;
cosLookup[15375] <= 0.096496303;
cosLookup[15376] <= 0.09640087;
cosLookup[15377] <= 0.096305436;
cosLookup[15378] <= 0.096210002;
cosLookup[15379] <= 0.096114567;
cosLookup[15380] <= 0.096019131;
cosLookup[15381] <= 0.095923693;
cosLookup[15382] <= 0.095828255;
cosLookup[15383] <= 0.095732817;
cosLookup[15384] <= 0.095637377;
cosLookup[15385] <= 0.095541936;
cosLookup[15386] <= 0.095446495;
cosLookup[15387] <= 0.095351052;
cosLookup[15388] <= 0.095255609;
cosLookup[15389] <= 0.095160165;
cosLookup[15390] <= 0.09506472;
cosLookup[15391] <= 0.094969274;
cosLookup[15392] <= 0.094873828;
cosLookup[15393] <= 0.09477838;
cosLookup[15394] <= 0.094682931;
cosLookup[15395] <= 0.094587482;
cosLookup[15396] <= 0.094492032;
cosLookup[15397] <= 0.094396581;
cosLookup[15398] <= 0.094301129;
cosLookup[15399] <= 0.094205676;
cosLookup[15400] <= 0.094110222;
cosLookup[15401] <= 0.094014768;
cosLookup[15402] <= 0.093919312;
cosLookup[15403] <= 0.093823856;
cosLookup[15404] <= 0.093728399;
cosLookup[15405] <= 0.093632941;
cosLookup[15406] <= 0.093537482;
cosLookup[15407] <= 0.093442022;
cosLookup[15408] <= 0.093346562;
cosLookup[15409] <= 0.0932511;
cosLookup[15410] <= 0.093155638;
cosLookup[15411] <= 0.093060175;
cosLookup[15412] <= 0.092964711;
cosLookup[15413] <= 0.092869246;
cosLookup[15414] <= 0.09277378;
cosLookup[15415] <= 0.092678314;
cosLookup[15416] <= 0.092582846;
cosLookup[15417] <= 0.092487378;
cosLookup[15418] <= 0.092391909;
cosLookup[15419] <= 0.092296439;
cosLookup[15420] <= 0.092200968;
cosLookup[15421] <= 0.092105497;
cosLookup[15422] <= 0.092010024;
cosLookup[15423] <= 0.091914551;
cosLookup[15424] <= 0.091819076;
cosLookup[15425] <= 0.091723601;
cosLookup[15426] <= 0.091628126;
cosLookup[15427] <= 0.091532649;
cosLookup[15428] <= 0.091437171;
cosLookup[15429] <= 0.091341693;
cosLookup[15430] <= 0.091246214;
cosLookup[15431] <= 0.091150733;
cosLookup[15432] <= 0.091055253;
cosLookup[15433] <= 0.090959771;
cosLookup[15434] <= 0.090864288;
cosLookup[15435] <= 0.090768805;
cosLookup[15436] <= 0.09067332;
cosLookup[15437] <= 0.090577835;
cosLookup[15438] <= 0.090482349;
cosLookup[15439] <= 0.090386863;
cosLookup[15440] <= 0.090291375;
cosLookup[15441] <= 0.090195887;
cosLookup[15442] <= 0.090100397;
cosLookup[15443] <= 0.090004907;
cosLookup[15444] <= 0.089909416;
cosLookup[15445] <= 0.089813925;
cosLookup[15446] <= 0.089718432;
cosLookup[15447] <= 0.089622939;
cosLookup[15448] <= 0.089527444;
cosLookup[15449] <= 0.089431949;
cosLookup[15450] <= 0.089336453;
cosLookup[15451] <= 0.089240957;
cosLookup[15452] <= 0.089145459;
cosLookup[15453] <= 0.089049961;
cosLookup[15454] <= 0.088954462;
cosLookup[15455] <= 0.088858962;
cosLookup[15456] <= 0.088763461;
cosLookup[15457] <= 0.088667959;
cosLookup[15458] <= 0.088572457;
cosLookup[15459] <= 0.088476954;
cosLookup[15460] <= 0.08838145;
cosLookup[15461] <= 0.088285945;
cosLookup[15462] <= 0.088190439;
cosLookup[15463] <= 0.088094933;
cosLookup[15464] <= 0.087999425;
cosLookup[15465] <= 0.087903917;
cosLookup[15466] <= 0.087808408;
cosLookup[15467] <= 0.087712899;
cosLookup[15468] <= 0.087617388;
cosLookup[15469] <= 0.087521877;
cosLookup[15470] <= 0.087426365;
cosLookup[15471] <= 0.087330852;
cosLookup[15472] <= 0.087235338;
cosLookup[15473] <= 0.087139824;
cosLookup[15474] <= 0.087044308;
cosLookup[15475] <= 0.086948792;
cosLookup[15476] <= 0.086853275;
cosLookup[15477] <= 0.086757757;
cosLookup[15478] <= 0.086662239;
cosLookup[15479] <= 0.08656672;
cosLookup[15480] <= 0.086471199;
cosLookup[15481] <= 0.086375679;
cosLookup[15482] <= 0.086280157;
cosLookup[15483] <= 0.086184634;
cosLookup[15484] <= 0.086089111;
cosLookup[15485] <= 0.085993587;
cosLookup[15486] <= 0.085898062;
cosLookup[15487] <= 0.085802536;
cosLookup[15488] <= 0.08570701;
cosLookup[15489] <= 0.085611483;
cosLookup[15490] <= 0.085515955;
cosLookup[15491] <= 0.085420426;
cosLookup[15492] <= 0.085324896;
cosLookup[15493] <= 0.085229366;
cosLookup[15494] <= 0.085133835;
cosLookup[15495] <= 0.085038303;
cosLookup[15496] <= 0.08494277;
cosLookup[15497] <= 0.084847237;
cosLookup[15498] <= 0.084751702;
cosLookup[15499] <= 0.084656167;
cosLookup[15500] <= 0.084560631;
cosLookup[15501] <= 0.084465095;
cosLookup[15502] <= 0.084369557;
cosLookup[15503] <= 0.084274019;
cosLookup[15504] <= 0.08417848;
cosLookup[15505] <= 0.08408294;
cosLookup[15506] <= 0.0839874;
cosLookup[15507] <= 0.083891859;
cosLookup[15508] <= 0.083796317;
cosLookup[15509] <= 0.083700774;
cosLookup[15510] <= 0.08360523;
cosLookup[15511] <= 0.083509686;
cosLookup[15512] <= 0.083414141;
cosLookup[15513] <= 0.083318595;
cosLookup[15514] <= 0.083223048;
cosLookup[15515] <= 0.083127501;
cosLookup[15516] <= 0.083031952;
cosLookup[15517] <= 0.082936404;
cosLookup[15518] <= 0.082840854;
cosLookup[15519] <= 0.082745303;
cosLookup[15520] <= 0.082649752;
cosLookup[15521] <= 0.0825542;
cosLookup[15522] <= 0.082458647;
cosLookup[15523] <= 0.082363094;
cosLookup[15524] <= 0.08226754;
cosLookup[15525] <= 0.082171985;
cosLookup[15526] <= 0.082076429;
cosLookup[15527] <= 0.081980872;
cosLookup[15528] <= 0.081885315;
cosLookup[15529] <= 0.081789757;
cosLookup[15530] <= 0.081694198;
cosLookup[15531] <= 0.081598639;
cosLookup[15532] <= 0.081503078;
cosLookup[15533] <= 0.081407517;
cosLookup[15534] <= 0.081311955;
cosLookup[15535] <= 0.081216393;
cosLookup[15536] <= 0.08112083;
cosLookup[15537] <= 0.081025266;
cosLookup[15538] <= 0.080929701;
cosLookup[15539] <= 0.080834135;
cosLookup[15540] <= 0.080738569;
cosLookup[15541] <= 0.080643002;
cosLookup[15542] <= 0.080547434;
cosLookup[15543] <= 0.080451866;
cosLookup[15544] <= 0.080356297;
cosLookup[15545] <= 0.080260727;
cosLookup[15546] <= 0.080165156;
cosLookup[15547] <= 0.080069584;
cosLookup[15548] <= 0.079974012;
cosLookup[15549] <= 0.079878439;
cosLookup[15550] <= 0.079782866;
cosLookup[15551] <= 0.079687291;
cosLookup[15552] <= 0.079591716;
cosLookup[15553] <= 0.07949614;
cosLookup[15554] <= 0.079400564;
cosLookup[15555] <= 0.079304987;
cosLookup[15556] <= 0.079209409;
cosLookup[15557] <= 0.07911383;
cosLookup[15558] <= 0.07901825;
cosLookup[15559] <= 0.07892267;
cosLookup[15560] <= 0.078827089;
cosLookup[15561] <= 0.078731507;
cosLookup[15562] <= 0.078635925;
cosLookup[15563] <= 0.078540342;
cosLookup[15564] <= 0.078444758;
cosLookup[15565] <= 0.078349174;
cosLookup[15566] <= 0.078253588;
cosLookup[15567] <= 0.078158002;
cosLookup[15568] <= 0.078062416;
cosLookup[15569] <= 0.077966828;
cosLookup[15570] <= 0.07787124;
cosLookup[15571] <= 0.077775651;
cosLookup[15572] <= 0.077680062;
cosLookup[15573] <= 0.077584471;
cosLookup[15574] <= 0.07748888;
cosLookup[15575] <= 0.077393289;
cosLookup[15576] <= 0.077297696;
cosLookup[15577] <= 0.077202103;
cosLookup[15578] <= 0.077106509;
cosLookup[15579] <= 0.077010915;
cosLookup[15580] <= 0.076915319;
cosLookup[15581] <= 0.076819723;
cosLookup[15582] <= 0.076724127;
cosLookup[15583] <= 0.076628529;
cosLookup[15584] <= 0.076532931;
cosLookup[15585] <= 0.076437332;
cosLookup[15586] <= 0.076341733;
cosLookup[15587] <= 0.076246133;
cosLookup[15588] <= 0.076150532;
cosLookup[15589] <= 0.07605493;
cosLookup[15590] <= 0.075959328;
cosLookup[15591] <= 0.075863725;
cosLookup[15592] <= 0.075768121;
cosLookup[15593] <= 0.075672517;
cosLookup[15594] <= 0.075576912;
cosLookup[15595] <= 0.075481306;
cosLookup[15596] <= 0.075385699;
cosLookup[15597] <= 0.075290092;
cosLookup[15598] <= 0.075194484;
cosLookup[15599] <= 0.075098876;
cosLookup[15600] <= 0.075003267;
cosLookup[15601] <= 0.074907657;
cosLookup[15602] <= 0.074812046;
cosLookup[15603] <= 0.074716435;
cosLookup[15604] <= 0.074620823;
cosLookup[15605] <= 0.07452521;
cosLookup[15606] <= 0.074429597;
cosLookup[15607] <= 0.074333983;
cosLookup[15608] <= 0.074238368;
cosLookup[15609] <= 0.074142753;
cosLookup[15610] <= 0.074047136;
cosLookup[15611] <= 0.07395152;
cosLookup[15612] <= 0.073855902;
cosLookup[15613] <= 0.073760284;
cosLookup[15614] <= 0.073664665;
cosLookup[15615] <= 0.073569046;
cosLookup[15616] <= 0.073473426;
cosLookup[15617] <= 0.073377805;
cosLookup[15618] <= 0.073282183;
cosLookup[15619] <= 0.073186561;
cosLookup[15620] <= 0.073090938;
cosLookup[15621] <= 0.072995315;
cosLookup[15622] <= 0.07289969;
cosLookup[15623] <= 0.072804066;
cosLookup[15624] <= 0.07270844;
cosLookup[15625] <= 0.072612814;
cosLookup[15626] <= 0.072517187;
cosLookup[15627] <= 0.072421559;
cosLookup[15628] <= 0.072325931;
cosLookup[15629] <= 0.072230302;
cosLookup[15630] <= 0.072134673;
cosLookup[15631] <= 0.072039043;
cosLookup[15632] <= 0.071943412;
cosLookup[15633] <= 0.07184778;
cosLookup[15634] <= 0.071752148;
cosLookup[15635] <= 0.071656515;
cosLookup[15636] <= 0.071560882;
cosLookup[15637] <= 0.071465247;
cosLookup[15638] <= 0.071369613;
cosLookup[15639] <= 0.071273977;
cosLookup[15640] <= 0.071178341;
cosLookup[15641] <= 0.071082704;
cosLookup[15642] <= 0.070987067;
cosLookup[15643] <= 0.070891429;
cosLookup[15644] <= 0.07079579;
cosLookup[15645] <= 0.070700151;
cosLookup[15646] <= 0.07060451;
cosLookup[15647] <= 0.07050887;
cosLookup[15648] <= 0.070413228;
cosLookup[15649] <= 0.070317586;
cosLookup[15650] <= 0.070221944;
cosLookup[15651] <= 0.070126301;
cosLookup[15652] <= 0.070030657;
cosLookup[15653] <= 0.069935012;
cosLookup[15654] <= 0.069839367;
cosLookup[15655] <= 0.069743721;
cosLookup[15656] <= 0.069648074;
cosLookup[15657] <= 0.069552427;
cosLookup[15658] <= 0.06945678;
cosLookup[15659] <= 0.069361131;
cosLookup[15660] <= 0.069265482;
cosLookup[15661] <= 0.069169832;
cosLookup[15662] <= 0.069074182;
cosLookup[15663] <= 0.068978531;
cosLookup[15664] <= 0.068882879;
cosLookup[15665] <= 0.068787227;
cosLookup[15666] <= 0.068691574;
cosLookup[15667] <= 0.068595921;
cosLookup[15668] <= 0.068500267;
cosLookup[15669] <= 0.068404612;
cosLookup[15670] <= 0.068308957;
cosLookup[15671] <= 0.068213301;
cosLookup[15672] <= 0.068117644;
cosLookup[15673] <= 0.068021987;
cosLookup[15674] <= 0.067926329;
cosLookup[15675] <= 0.06783067;
cosLookup[15676] <= 0.067735011;
cosLookup[15677] <= 0.067639351;
cosLookup[15678] <= 0.067543691;
cosLookup[15679] <= 0.06744803;
cosLookup[15680] <= 0.067352368;
cosLookup[15681] <= 0.067256706;
cosLookup[15682] <= 0.067161043;
cosLookup[15683] <= 0.06706538;
cosLookup[15684] <= 0.066969716;
cosLookup[15685] <= 0.066874051;
cosLookup[15686] <= 0.066778386;
cosLookup[15687] <= 0.06668272;
cosLookup[15688] <= 0.066587053;
cosLookup[15689] <= 0.066491386;
cosLookup[15690] <= 0.066395718;
cosLookup[15691] <= 0.06630005;
cosLookup[15692] <= 0.066204381;
cosLookup[15693] <= 0.066108711;
cosLookup[15694] <= 0.066013041;
cosLookup[15695] <= 0.06591737;
cosLookup[15696] <= 0.065821699;
cosLookup[15697] <= 0.065726027;
cosLookup[15698] <= 0.065630354;
cosLookup[15699] <= 0.065534681;
cosLookup[15700] <= 0.065439007;
cosLookup[15701] <= 0.065343333;
cosLookup[15702] <= 0.065247658;
cosLookup[15703] <= 0.065151982;
cosLookup[15704] <= 0.065056306;
cosLookup[15705] <= 0.064960629;
cosLookup[15706] <= 0.064864951;
cosLookup[15707] <= 0.064769273;
cosLookup[15708] <= 0.064673595;
cosLookup[15709] <= 0.064577916;
cosLookup[15710] <= 0.064482236;
cosLookup[15711] <= 0.064386555;
cosLookup[15712] <= 0.064290874;
cosLookup[15713] <= 0.064195193;
cosLookup[15714] <= 0.064099511;
cosLookup[15715] <= 0.064003828;
cosLookup[15716] <= 0.063908144;
cosLookup[15717] <= 0.06381246;
cosLookup[15718] <= 0.063716776;
cosLookup[15719] <= 0.063621091;
cosLookup[15720] <= 0.063525405;
cosLookup[15721] <= 0.063429719;
cosLookup[15722] <= 0.063334032;
cosLookup[15723] <= 0.063238345;
cosLookup[15724] <= 0.063142656;
cosLookup[15725] <= 0.063046968;
cosLookup[15726] <= 0.062951279;
cosLookup[15727] <= 0.062855589;
cosLookup[15728] <= 0.062759899;
cosLookup[15729] <= 0.062664208;
cosLookup[15730] <= 0.062568516;
cosLookup[15731] <= 0.062472824;
cosLookup[15732] <= 0.062377131;
cosLookup[15733] <= 0.062281438;
cosLookup[15734] <= 0.062185744;
cosLookup[15735] <= 0.06209005;
cosLookup[15736] <= 0.061994355;
cosLookup[15737] <= 0.06189866;
cosLookup[15738] <= 0.061802963;
cosLookup[15739] <= 0.061707267;
cosLookup[15740] <= 0.06161157;
cosLookup[15741] <= 0.061515872;
cosLookup[15742] <= 0.061420173;
cosLookup[15743] <= 0.061324475;
cosLookup[15744] <= 0.061228775;
cosLookup[15745] <= 0.061133075;
cosLookup[15746] <= 0.061037374;
cosLookup[15747] <= 0.060941673;
cosLookup[15748] <= 0.060845972;
cosLookup[15749] <= 0.060750269;
cosLookup[15750] <= 0.060654566;
cosLookup[15751] <= 0.060558863;
cosLookup[15752] <= 0.060463159;
cosLookup[15753] <= 0.060367455;
cosLookup[15754] <= 0.06027175;
cosLookup[15755] <= 0.060176044;
cosLookup[15756] <= 0.060080338;
cosLookup[15757] <= 0.059984631;
cosLookup[15758] <= 0.059888924;
cosLookup[15759] <= 0.059793216;
cosLookup[15760] <= 0.059697508;
cosLookup[15761] <= 0.059601799;
cosLookup[15762] <= 0.059506089;
cosLookup[15763] <= 0.059410379;
cosLookup[15764] <= 0.059314669;
cosLookup[15765] <= 0.059218957;
cosLookup[15766] <= 0.059123246;
cosLookup[15767] <= 0.059027534;
cosLookup[15768] <= 0.058931821;
cosLookup[15769] <= 0.058836108;
cosLookup[15770] <= 0.058740394;
cosLookup[15771] <= 0.058644679;
cosLookup[15772] <= 0.058548964;
cosLookup[15773] <= 0.058453249;
cosLookup[15774] <= 0.058357533;
cosLookup[15775] <= 0.058261816;
cosLookup[15776] <= 0.058166099;
cosLookup[15777] <= 0.058070382;
cosLookup[15778] <= 0.057974664;
cosLookup[15779] <= 0.057878945;
cosLookup[15780] <= 0.057783226;
cosLookup[15781] <= 0.057687506;
cosLookup[15782] <= 0.057591786;
cosLookup[15783] <= 0.057496065;
cosLookup[15784] <= 0.057400344;
cosLookup[15785] <= 0.057304622;
cosLookup[15786] <= 0.0572089;
cosLookup[15787] <= 0.057113177;
cosLookup[15788] <= 0.057017453;
cosLookup[15789] <= 0.056921729;
cosLookup[15790] <= 0.056826005;
cosLookup[15791] <= 0.05673028;
cosLookup[15792] <= 0.056634554;
cosLookup[15793] <= 0.056538828;
cosLookup[15794] <= 0.056443102;
cosLookup[15795] <= 0.056347375;
cosLookup[15796] <= 0.056251647;
cosLookup[15797] <= 0.056155919;
cosLookup[15798] <= 0.056060191;
cosLookup[15799] <= 0.055964461;
cosLookup[15800] <= 0.055868732;
cosLookup[15801] <= 0.055773002;
cosLookup[15802] <= 0.055677271;
cosLookup[15803] <= 0.05558154;
cosLookup[15804] <= 0.055485808;
cosLookup[15805] <= 0.055390076;
cosLookup[15806] <= 0.055294343;
cosLookup[15807] <= 0.05519861;
cosLookup[15808] <= 0.055102876;
cosLookup[15809] <= 0.055007142;
cosLookup[15810] <= 0.054911407;
cosLookup[15811] <= 0.054815672;
cosLookup[15812] <= 0.054719936;
cosLookup[15813] <= 0.0546242;
cosLookup[15814] <= 0.054528463;
cosLookup[15815] <= 0.054432726;
cosLookup[15816] <= 0.054336988;
cosLookup[15817] <= 0.05424125;
cosLookup[15818] <= 0.054145511;
cosLookup[15819] <= 0.054049772;
cosLookup[15820] <= 0.053954032;
cosLookup[15821] <= 0.053858292;
cosLookup[15822] <= 0.053762551;
cosLookup[15823] <= 0.05366681;
cosLookup[15824] <= 0.053571068;
cosLookup[15825] <= 0.053475326;
cosLookup[15826] <= 0.053379583;
cosLookup[15827] <= 0.05328384;
cosLookup[15828] <= 0.053188097;
cosLookup[15829] <= 0.053092352;
cosLookup[15830] <= 0.052996608;
cosLookup[15831] <= 0.052900863;
cosLookup[15832] <= 0.052805117;
cosLookup[15833] <= 0.052709371;
cosLookup[15834] <= 0.052613624;
cosLookup[15835] <= 0.052517877;
cosLookup[15836] <= 0.052422129;
cosLookup[15837] <= 0.052326381;
cosLookup[15838] <= 0.052230633;
cosLookup[15839] <= 0.052134884;
cosLookup[15840] <= 0.052039134;
cosLookup[15841] <= 0.051943384;
cosLookup[15842] <= 0.051847634;
cosLookup[15843] <= 0.051751883;
cosLookup[15844] <= 0.051656132;
cosLookup[15845] <= 0.05156038;
cosLookup[15846] <= 0.051464627;
cosLookup[15847] <= 0.051368875;
cosLookup[15848] <= 0.051273121;
cosLookup[15849] <= 0.051177367;
cosLookup[15850] <= 0.051081613;
cosLookup[15851] <= 0.050985858;
cosLookup[15852] <= 0.050890103;
cosLookup[15853] <= 0.050794348;
cosLookup[15854] <= 0.050698592;
cosLookup[15855] <= 0.050602835;
cosLookup[15856] <= 0.050507078;
cosLookup[15857] <= 0.05041132;
cosLookup[15858] <= 0.050315562;
cosLookup[15859] <= 0.050219804;
cosLookup[15860] <= 0.050124045;
cosLookup[15861] <= 0.050028286;
cosLookup[15862] <= 0.049932526;
cosLookup[15863] <= 0.049836766;
cosLookup[15864] <= 0.049741005;
cosLookup[15865] <= 0.049645244;
cosLookup[15866] <= 0.049549482;
cosLookup[15867] <= 0.04945372;
cosLookup[15868] <= 0.049357957;
cosLookup[15869] <= 0.049262194;
cosLookup[15870] <= 0.049166431;
cosLookup[15871] <= 0.049070667;
cosLookup[15872] <= 0.048974903;
cosLookup[15873] <= 0.048879138;
cosLookup[15874] <= 0.048783372;
cosLookup[15875] <= 0.048687607;
cosLookup[15876] <= 0.048591841;
cosLookup[15877] <= 0.048496074;
cosLookup[15878] <= 0.048400307;
cosLookup[15879] <= 0.048304539;
cosLookup[15880] <= 0.048208771;
cosLookup[15881] <= 0.048113003;
cosLookup[15882] <= 0.048017234;
cosLookup[15883] <= 0.047921465;
cosLookup[15884] <= 0.047825695;
cosLookup[15885] <= 0.047729925;
cosLookup[15886] <= 0.047634155;
cosLookup[15887] <= 0.047538383;
cosLookup[15888] <= 0.047442612;
cosLookup[15889] <= 0.04734684;
cosLookup[15890] <= 0.047251068;
cosLookup[15891] <= 0.047155295;
cosLookup[15892] <= 0.047059522;
cosLookup[15893] <= 0.046963748;
cosLookup[15894] <= 0.046867974;
cosLookup[15895] <= 0.0467722;
cosLookup[15896] <= 0.046676425;
cosLookup[15897] <= 0.046580649;
cosLookup[15898] <= 0.046484873;
cosLookup[15899] <= 0.046389097;
cosLookup[15900] <= 0.046293321;
cosLookup[15901] <= 0.046197544;
cosLookup[15902] <= 0.046101766;
cosLookup[15903] <= 0.046005988;
cosLookup[15904] <= 0.04591021;
cosLookup[15905] <= 0.045814431;
cosLookup[15906] <= 0.045718652;
cosLookup[15907] <= 0.045622872;
cosLookup[15908] <= 0.045527092;
cosLookup[15909] <= 0.045431312;
cosLookup[15910] <= 0.045335531;
cosLookup[15911] <= 0.04523975;
cosLookup[15912] <= 0.045143968;
cosLookup[15913] <= 0.045048186;
cosLookup[15914] <= 0.044952403;
cosLookup[15915] <= 0.04485662;
cosLookup[15916] <= 0.044760837;
cosLookup[15917] <= 0.044665053;
cosLookup[15918] <= 0.044569269;
cosLookup[15919] <= 0.044473485;
cosLookup[15920] <= 0.0443777;
cosLookup[15921] <= 0.044281914;
cosLookup[15922] <= 0.044186128;
cosLookup[15923] <= 0.044090342;
cosLookup[15924] <= 0.043994555;
cosLookup[15925] <= 0.043898768;
cosLookup[15926] <= 0.043802981;
cosLookup[15927] <= 0.043707193;
cosLookup[15928] <= 0.043611405;
cosLookup[15929] <= 0.043515616;
cosLookup[15930] <= 0.043419827;
cosLookup[15931] <= 0.043324038;
cosLookup[15932] <= 0.043228248;
cosLookup[15933] <= 0.043132458;
cosLookup[15934] <= 0.043036667;
cosLookup[15935] <= 0.042940876;
cosLookup[15936] <= 0.042845085;
cosLookup[15937] <= 0.042749293;
cosLookup[15938] <= 0.042653501;
cosLookup[15939] <= 0.042557708;
cosLookup[15940] <= 0.042461915;
cosLookup[15941] <= 0.042366122;
cosLookup[15942] <= 0.042270328;
cosLookup[15943] <= 0.042174534;
cosLookup[15944] <= 0.042078739;
cosLookup[15945] <= 0.041982945;
cosLookup[15946] <= 0.041887149;
cosLookup[15947] <= 0.041791353;
cosLookup[15948] <= 0.041695557;
cosLookup[15949] <= 0.041599761;
cosLookup[15950] <= 0.041503964;
cosLookup[15951] <= 0.041408167;
cosLookup[15952] <= 0.041312369;
cosLookup[15953] <= 0.041216571;
cosLookup[15954] <= 0.041120773;
cosLookup[15955] <= 0.041024974;
cosLookup[15956] <= 0.040929175;
cosLookup[15957] <= 0.040833376;
cosLookup[15958] <= 0.040737576;
cosLookup[15959] <= 0.040641775;
cosLookup[15960] <= 0.040545975;
cosLookup[15961] <= 0.040450174;
cosLookup[15962] <= 0.040354372;
cosLookup[15963] <= 0.040258571;
cosLookup[15964] <= 0.040162769;
cosLookup[15965] <= 0.040066966;
cosLookup[15966] <= 0.039971163;
cosLookup[15967] <= 0.03987536;
cosLookup[15968] <= 0.039779557;
cosLookup[15969] <= 0.039683753;
cosLookup[15970] <= 0.039587948;
cosLookup[15971] <= 0.039492144;
cosLookup[15972] <= 0.039396339;
cosLookup[15973] <= 0.039300533;
cosLookup[15974] <= 0.039204727;
cosLookup[15975] <= 0.039108921;
cosLookup[15976] <= 0.039013115;
cosLookup[15977] <= 0.038917308;
cosLookup[15978] <= 0.038821501;
cosLookup[15979] <= 0.038725693;
cosLookup[15980] <= 0.038629885;
cosLookup[15981] <= 0.038534077;
cosLookup[15982] <= 0.038438268;
cosLookup[15983] <= 0.038342459;
cosLookup[15984] <= 0.03824665;
cosLookup[15985] <= 0.03815084;
cosLookup[15986] <= 0.03805503;
cosLookup[15987] <= 0.03795922;
cosLookup[15988] <= 0.037863409;
cosLookup[15989] <= 0.037767598;
cosLookup[15990] <= 0.037671787;
cosLookup[15991] <= 0.037575975;
cosLookup[15992] <= 0.037480163;
cosLookup[15993] <= 0.037384351;
cosLookup[15994] <= 0.037288538;
cosLookup[15995] <= 0.037192725;
cosLookup[15996] <= 0.037096911;
cosLookup[15997] <= 0.037001097;
cosLookup[15998] <= 0.036905283;
cosLookup[15999] <= 0.036809469;
cosLookup[16000] <= 0.036713654;
cosLookup[16001] <= 0.036617839;
cosLookup[16002] <= 0.036522023;
cosLookup[16003] <= 0.036426207;
cosLookup[16004] <= 0.036330391;
cosLookup[16005] <= 0.036234574;
cosLookup[16006] <= 0.036138758;
cosLookup[16007] <= 0.03604294;
cosLookup[16008] <= 0.035947123;
cosLookup[16009] <= 0.035851305;
cosLookup[16010] <= 0.035755487;
cosLookup[16011] <= 0.035659668;
cosLookup[16012] <= 0.03556385;
cosLookup[16013] <= 0.03546803;
cosLookup[16014] <= 0.035372211;
cosLookup[16015] <= 0.035276391;
cosLookup[16016] <= 0.035180571;
cosLookup[16017] <= 0.035084751;
cosLookup[16018] <= 0.03498893;
cosLookup[16019] <= 0.034893109;
cosLookup[16020] <= 0.034797287;
cosLookup[16021] <= 0.034701465;
cosLookup[16022] <= 0.034605643;
cosLookup[16023] <= 0.034509821;
cosLookup[16024] <= 0.034413998;
cosLookup[16025] <= 0.034318175;
cosLookup[16026] <= 0.034222352;
cosLookup[16027] <= 0.034126528;
cosLookup[16028] <= 0.034030704;
cosLookup[16029] <= 0.03393488;
cosLookup[16030] <= 0.033839055;
cosLookup[16031] <= 0.033743231;
cosLookup[16032] <= 0.033647405;
cosLookup[16033] <= 0.03355158;
cosLookup[16034] <= 0.033455754;
cosLookup[16035] <= 0.033359928;
cosLookup[16036] <= 0.033264101;
cosLookup[16037] <= 0.033168275;
cosLookup[16038] <= 0.033072448;
cosLookup[16039] <= 0.03297662;
cosLookup[16040] <= 0.032880793;
cosLookup[16041] <= 0.032784965;
cosLookup[16042] <= 0.032689136;
cosLookup[16043] <= 0.032593308;
cosLookup[16044] <= 0.032497479;
cosLookup[16045] <= 0.03240165;
cosLookup[16046] <= 0.03230582;
cosLookup[16047] <= 0.032209991;
cosLookup[16048] <= 0.032114161;
cosLookup[16049] <= 0.03201833;
cosLookup[16050] <= 0.0319225;
cosLookup[16051] <= 0.031826669;
cosLookup[16052] <= 0.031730837;
cosLookup[16053] <= 0.031635006;
cosLookup[16054] <= 0.031539174;
cosLookup[16055] <= 0.031443342;
cosLookup[16056] <= 0.03134751;
cosLookup[16057] <= 0.031251677;
cosLookup[16058] <= 0.031155844;
cosLookup[16059] <= 0.031060011;
cosLookup[16060] <= 0.030964177;
cosLookup[16061] <= 0.030868343;
cosLookup[16062] <= 0.030772509;
cosLookup[16063] <= 0.030676675;
cosLookup[16064] <= 0.03058084;
cosLookup[16065] <= 0.030485005;
cosLookup[16066] <= 0.03038917;
cosLookup[16067] <= 0.030293335;
cosLookup[16068] <= 0.030197499;
cosLookup[16069] <= 0.030101663;
cosLookup[16070] <= 0.030005826;
cosLookup[16071] <= 0.02990999;
cosLookup[16072] <= 0.029814153;
cosLookup[16073] <= 0.029718316;
cosLookup[16074] <= 0.029622478;
cosLookup[16075] <= 0.029526641;
cosLookup[16076] <= 0.029430803;
cosLookup[16077] <= 0.029334964;
cosLookup[16078] <= 0.029239126;
cosLookup[16079] <= 0.029143287;
cosLookup[16080] <= 0.029047448;
cosLookup[16081] <= 0.028951609;
cosLookup[16082] <= 0.028855769;
cosLookup[16083] <= 0.028759929;
cosLookup[16084] <= 0.028664089;
cosLookup[16085] <= 0.028568249;
cosLookup[16086] <= 0.028472408;
cosLookup[16087] <= 0.028376567;
cosLookup[16088] <= 0.028280726;
cosLookup[16089] <= 0.028184885;
cosLookup[16090] <= 0.028089043;
cosLookup[16091] <= 0.027993201;
cosLookup[16092] <= 0.027897359;
cosLookup[16093] <= 0.027801516;
cosLookup[16094] <= 0.027705673;
cosLookup[16095] <= 0.027609831;
cosLookup[16096] <= 0.027513987;
cosLookup[16097] <= 0.027418144;
cosLookup[16098] <= 0.0273223;
cosLookup[16099] <= 0.027226456;
cosLookup[16100] <= 0.027130612;
cosLookup[16101] <= 0.027034767;
cosLookup[16102] <= 0.026938923;
cosLookup[16103] <= 0.026843078;
cosLookup[16104] <= 0.026747232;
cosLookup[16105] <= 0.026651387;
cosLookup[16106] <= 0.026555541;
cosLookup[16107] <= 0.026459695;
cosLookup[16108] <= 0.026363849;
cosLookup[16109] <= 0.026268003;
cosLookup[16110] <= 0.026172156;
cosLookup[16111] <= 0.026076309;
cosLookup[16112] <= 0.025980462;
cosLookup[16113] <= 0.025884614;
cosLookup[16114] <= 0.025788767;
cosLookup[16115] <= 0.025692919;
cosLookup[16116] <= 0.025597071;
cosLookup[16117] <= 0.025501222;
cosLookup[16118] <= 0.025405374;
cosLookup[16119] <= 0.025309525;
cosLookup[16120] <= 0.025213676;
cosLookup[16121] <= 0.025117827;
cosLookup[16122] <= 0.025021977;
cosLookup[16123] <= 0.024926127;
cosLookup[16124] <= 0.024830277;
cosLookup[16125] <= 0.024734427;
cosLookup[16126] <= 0.024638577;
cosLookup[16127] <= 0.024542726;
cosLookup[16128] <= 0.024446875;
cosLookup[16129] <= 0.024351024;
cosLookup[16130] <= 0.024255173;
cosLookup[16131] <= 0.024159321;
cosLookup[16132] <= 0.02406347;
cosLookup[16133] <= 0.023967618;
cosLookup[16134] <= 0.023871765;
cosLookup[16135] <= 0.023775913;
cosLookup[16136] <= 0.02368006;
cosLookup[16137] <= 0.023584207;
cosLookup[16138] <= 0.023488354;
cosLookup[16139] <= 0.023392501;
cosLookup[16140] <= 0.023296647;
cosLookup[16141] <= 0.023200794;
cosLookup[16142] <= 0.02310494;
cosLookup[16143] <= 0.023009086;
cosLookup[16144] <= 0.022913231;
cosLookup[16145] <= 0.022817377;
cosLookup[16146] <= 0.022721522;
cosLookup[16147] <= 0.022625667;
cosLookup[16148] <= 0.022529812;
cosLookup[16149] <= 0.022433956;
cosLookup[16150] <= 0.022338101;
cosLookup[16151] <= 0.022242245;
cosLookup[16152] <= 0.022146389;
cosLookup[16153] <= 0.022050532;
cosLookup[16154] <= 0.021954676;
cosLookup[16155] <= 0.021858819;
cosLookup[16156] <= 0.021762963;
cosLookup[16157] <= 0.021667106;
cosLookup[16158] <= 0.021571248;
cosLookup[16159] <= 0.021475391;
cosLookup[16160] <= 0.021379533;
cosLookup[16161] <= 0.021283675;
cosLookup[16162] <= 0.021187817;
cosLookup[16163] <= 0.021091959;
cosLookup[16164] <= 0.020996101;
cosLookup[16165] <= 0.020900242;
cosLookup[16166] <= 0.020804383;
cosLookup[16167] <= 0.020708524;
cosLookup[16168] <= 0.020612665;
cosLookup[16169] <= 0.020516806;
cosLookup[16170] <= 0.020420946;
cosLookup[16171] <= 0.020325086;
cosLookup[16172] <= 0.020229226;
cosLookup[16173] <= 0.020133366;
cosLookup[16174] <= 0.020037506;
cosLookup[16175] <= 0.019941646;
cosLookup[16176] <= 0.019845785;
cosLookup[16177] <= 0.019749924;
cosLookup[16178] <= 0.019654063;
cosLookup[16179] <= 0.019558202;
cosLookup[16180] <= 0.01946234;
cosLookup[16181] <= 0.019366479;
cosLookup[16182] <= 0.019270617;
cosLookup[16183] <= 0.019174755;
cosLookup[16184] <= 0.019078893;
cosLookup[16185] <= 0.018983031;
cosLookup[16186] <= 0.018887168;
cosLookup[16187] <= 0.018791306;
cosLookup[16188] <= 0.018695443;
cosLookup[16189] <= 0.01859958;
cosLookup[16190] <= 0.018503717;
cosLookup[16191] <= 0.018407853;
cosLookup[16192] <= 0.01831199;
cosLookup[16193] <= 0.018216126;
cosLookup[16194] <= 0.018120262;
cosLookup[16195] <= 0.018024398;
cosLookup[16196] <= 0.017928534;
cosLookup[16197] <= 0.01783267;
cosLookup[16198] <= 0.017736805;
cosLookup[16199] <= 0.017640941;
cosLookup[16200] <= 0.017545076;
cosLookup[16201] <= 0.017449211;
cosLookup[16202] <= 0.017353346;
cosLookup[16203] <= 0.017257481;
cosLookup[16204] <= 0.017161615;
cosLookup[16205] <= 0.017065749;
cosLookup[16206] <= 0.016969884;
cosLookup[16207] <= 0.016874018;
cosLookup[16208] <= 0.016778152;
cosLookup[16209] <= 0.016682285;
cosLookup[16210] <= 0.016586419;
cosLookup[16211] <= 0.016490553;
cosLookup[16212] <= 0.016394686;
cosLookup[16213] <= 0.016298819;
cosLookup[16214] <= 0.016202952;
cosLookup[16215] <= 0.016107085;
cosLookup[16216] <= 0.016011218;
cosLookup[16217] <= 0.01591535;
cosLookup[16218] <= 0.015819483;
cosLookup[16219] <= 0.015723615;
cosLookup[16220] <= 0.015627747;
cosLookup[16221] <= 0.015531879;
cosLookup[16222] <= 0.015436011;
cosLookup[16223] <= 0.015340142;
cosLookup[16224] <= 0.015244274;
cosLookup[16225] <= 0.015148405;
cosLookup[16226] <= 0.015052537;
cosLookup[16227] <= 0.014956668;
cosLookup[16228] <= 0.014860799;
cosLookup[16229] <= 0.01476493;
cosLookup[16230] <= 0.014669061;
cosLookup[16231] <= 0.014573191;
cosLookup[16232] <= 0.014477322;
cosLookup[16233] <= 0.014381452;
cosLookup[16234] <= 0.014285582;
cosLookup[16235] <= 0.014189712;
cosLookup[16236] <= 0.014093842;
cosLookup[16237] <= 0.013997972;
cosLookup[16238] <= 0.013902102;
cosLookup[16239] <= 0.013806231;
cosLookup[16240] <= 0.013710361;
cosLookup[16241] <= 0.01361449;
cosLookup[16242] <= 0.013518619;
cosLookup[16243] <= 0.013422748;
cosLookup[16244] <= 0.013326877;
cosLookup[16245] <= 0.013231006;
cosLookup[16246] <= 0.013135134;
cosLookup[16247] <= 0.013039263;
cosLookup[16248] <= 0.012943391;
cosLookup[16249] <= 0.01284752;
cosLookup[16250] <= 0.012751648;
cosLookup[16251] <= 0.012655776;
cosLookup[16252] <= 0.012559904;
cosLookup[16253] <= 0.012464032;
cosLookup[16254] <= 0.01236816;
cosLookup[16255] <= 0.012272287;
cosLookup[16256] <= 0.012176415;
cosLookup[16257] <= 0.012080542;
cosLookup[16258] <= 0.011984669;
cosLookup[16259] <= 0.011888797;
cosLookup[16260] <= 0.011792924;
cosLookup[16261] <= 0.011697051;
cosLookup[16262] <= 0.011601178;
cosLookup[16263] <= 0.011505304;
cosLookup[16264] <= 0.011409431;
cosLookup[16265] <= 0.011313557;
cosLookup[16266] <= 0.011217684;
cosLookup[16267] <= 0.01112181;
cosLookup[16268] <= 0.011025936;
cosLookup[16269] <= 0.010930063;
cosLookup[16270] <= 0.010834189;
cosLookup[16271] <= 0.010738315;
cosLookup[16272] <= 0.01064244;
cosLookup[16273] <= 0.010546566;
cosLookup[16274] <= 0.010450692;
cosLookup[16275] <= 0.010354817;
cosLookup[16276] <= 0.010258943;
cosLookup[16277] <= 0.010163068;
cosLookup[16278] <= 0.010067193;
cosLookup[16279] <= 0.009971318;
cosLookup[16280] <= 0.009875444;
cosLookup[16281] <= 0.009779569;
cosLookup[16282] <= 0.009683693;
cosLookup[16283] <= 0.009587818;
cosLookup[16284] <= 0.009491943;
cosLookup[16285] <= 0.009396068;
cosLookup[16286] <= 0.009300192;
cosLookup[16287] <= 0.009204317;
cosLookup[16288] <= 0.009108441;
cosLookup[16289] <= 0.009012565;
cosLookup[16290] <= 0.008916689;
cosLookup[16291] <= 0.008820814;
cosLookup[16292] <= 0.008724938;
cosLookup[16293] <= 0.008629062;
cosLookup[16294] <= 0.008533185;
cosLookup[16295] <= 0.008437309;
cosLookup[16296] <= 0.008341433;
cosLookup[16297] <= 0.008245557;
cosLookup[16298] <= 0.00814968;
cosLookup[16299] <= 0.008053804;
cosLookup[16300] <= 0.007957927;
cosLookup[16301] <= 0.00786205;
cosLookup[16302] <= 0.007766174;
cosLookup[16303] <= 0.007670297;
cosLookup[16304] <= 0.00757442;
cosLookup[16305] <= 0.007478543;
cosLookup[16306] <= 0.007382666;
cosLookup[16307] <= 0.007286789;
cosLookup[16308] <= 0.007190912;
cosLookup[16309] <= 0.007095035;
cosLookup[16310] <= 0.006999157;
cosLookup[16311] <= 0.00690328;
cosLookup[16312] <= 0.006807403;
cosLookup[16313] <= 0.006711525;
cosLookup[16314] <= 0.006615648;
cosLookup[16315] <= 0.00651977;
cosLookup[16316] <= 0.006423892;
cosLookup[16317] <= 0.006328015;
cosLookup[16318] <= 0.006232137;
cosLookup[16319] <= 0.006136259;
cosLookup[16320] <= 0.006040381;
cosLookup[16321] <= 0.005944503;
cosLookup[16322] <= 0.005848625;
cosLookup[16323] <= 0.005752747;
cosLookup[16324] <= 0.005656869;
cosLookup[16325] <= 0.005560991;
cosLookup[16326] <= 0.005465113;
cosLookup[16327] <= 0.005369235;
cosLookup[16328] <= 0.005273356;
cosLookup[16329] <= 0.005177478;
cosLookup[16330] <= 0.0050816;
cosLookup[16331] <= 0.004985721;
cosLookup[16332] <= 0.004889843;
cosLookup[16333] <= 0.004793964;
cosLookup[16334] <= 0.004698086;
cosLookup[16335] <= 0.004602207;
cosLookup[16336] <= 0.004506328;
cosLookup[16337] <= 0.00441045;
cosLookup[16338] <= 0.004314571;
cosLookup[16339] <= 0.004218692;
cosLookup[16340] <= 0.004122813;
cosLookup[16341] <= 0.004026934;
cosLookup[16342] <= 0.003931056;
cosLookup[16343] <= 0.003835177;
cosLookup[16344] <= 0.003739298;
cosLookup[16345] <= 0.003643419;
cosLookup[16346] <= 0.00354754;
cosLookup[16347] <= 0.003451661;
cosLookup[16348] <= 0.003355781;
cosLookup[16349] <= 0.003259902;
cosLookup[16350] <= 0.003164023;
cosLookup[16351] <= 0.003068144;
cosLookup[16352] <= 0.002972265;
cosLookup[16353] <= 0.002876386;
cosLookup[16354] <= 0.002780506;
cosLookup[16355] <= 0.002684627;
cosLookup[16356] <= 0.002588748;
cosLookup[16357] <= 0.002492868;
cosLookup[16358] <= 0.002396989;
cosLookup[16359] <= 0.00230111;
cosLookup[16360] <= 0.00220523;
cosLookup[16361] <= 0.002109351;
cosLookup[16362] <= 0.002013471;
cosLookup[16363] <= 0.001917592;
cosLookup[16364] <= 0.001821712;
cosLookup[16365] <= 0.001725833;
cosLookup[16366] <= 0.001629953;
cosLookup[16367] <= 0.001534074;
cosLookup[16368] <= 0.001438194;
cosLookup[16369] <= 0.001342315;
cosLookup[16370] <= 0.001246435;
cosLookup[16371] <= 0.001150556;
cosLookup[16372] <= 0.001054676;
cosLookup[16373] <= 0.000958796;
cosLookup[16374] <= 0.000862917;
cosLookup[16375] <= 0.000767037;
cosLookup[16376] <= 0.000671158;
cosLookup[16377] <= 0.000575278;
cosLookup[16378] <= 0.000479398;
cosLookup[16379] <= 0.000383519;
cosLookup[16380] <= 0.000287639;
cosLookup[16381] <= 0.000191759;
cosLookup[16382] <= 0.0000958797;
cosLookup[16383] <= 6.12323E-17;
end

always @(x_sign)
begin
  if (x_sign == 1)
    assign g0 = -1*cosLookup[x_g_a];
  else
    assign g0 = cosLookup[x_g_a];
end

always @(y_sign)
begin
  if (y_sign == 1)
    assign g1 = -1*cosLookup[(1-2^-14) - x_g_a];
  else
    assign g1 = cosLookup[(1-2^-14) - x_g_a];
end

endmodule
